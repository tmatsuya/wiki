`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWuVD2G72UtjuvPh3IeG66mSo8uh/WEmRhJNlGQFER2voyHM6BgvOanMRJXtLg/2hJc5lS3PNilP
5zc0eSWvbw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GEiob5VmqGPB94ZQvO3SCyYhKMEhsy0Wwi7+oi28I+YKC7DjOHO3KcXgywz5q5Qh+dtSux1WpQYp
QZIHYrSpA7ceCJlnnG6Mv6631b2jfKunXY/u8J5KVsyhLv9BZ0fBOhw3iQbMPpnm72M8AoHj0lfG
sRTl49fEJ9sj4wUGE9Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ArpfjbVny9rahsVWoBweT7W/nHgi71tEonoV7bi6MH008LKUfazmWu+VAkWcNcoip795tzxWBL+K
xuyiY8Zbg3Gew46gUCQhAB8YLzqHlw1E0c9b2Xv8trOdVNZnNMEDvSqu9lTU+8ovaJXzJ+wkxhof
SwnNyR0tLmAyPQj8SM9JiHv37M0SHdOtOmNsYsLlx2OivNSXUOhUS08EyYy4blkopKTY+4GwG6Aj
EPhwCbaXB+/t1f1xpBT+2iRmSov0JoUiDgKU4YRARD4WreFKu3CVZMSlhMgalJVdGtE+yXUhChLJ
j/3pR8xc0NJtASb9KfW5ZK6sqI69z4uOIbqEsQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s7dFx2k3cHvygDkH+HoNU/iixuns48H18ck5fLM/YzjzgJb8uTWSv16RkFaFc9GXuI3UOarjVWsa
RaIDj9KdgGQQEXF8nBGTtZquli+JWdkGDv95zX8nxdnNHFqhkce7xA9ENDwUEAimiEWyX5BQbRjN
1nC30ar/it5plXYQEys=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IxxAx+cFNzqIiw/JjrHbXr5LH9yLe9OOXVZyHq45SCRFb3nXVUWnJMqFQ/2uwEyiLlv3zVUE+clq
kjNqmf6p7fE+MM14OSTGUBWFrCARbgzxuuPqJIYGsUqT2ysBcO28WhltXcHt0ijaVeE96Y+3vpfo
ibE/hNEi2efnsceXZNwx8qJu2prL+PrqLAIfuMI+eLcv9O7Ln1xQXx1CQpv9ZlwZ3eNWW1AG7j30
2kPZNPwJkpy6oW2aUY36sqzcJY95gv/4RDHDpP3HfSUhJ25QaenSQ1L5H539rTTk+M/WqePoJ4ME
FQ7dLrUIzlkfV1iHJ9GHmdqTJy/o2MHe3ujHyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12368)
`protect data_block
M3puya94M7ifbmnL3Y1DZBg20Fup9pAzDPE6Vy2Rm/Zj2GY0PBMjwHDZqIjHXyJZ+54/c2rGFEC8
Ki1ZqY2YN+/a6NiLwKtJOGc3VRDrslo/s7AUuntBBr64Qt7qxHJa8kmeXrVjWJFj+Zx+j5/KNeBG
9ai84upCrtwUEXOu7E4w3R//Qzcx542z1x/pQCZFQ1yovMeqVk3N3VUGbvJl+QiiqkPkwHK4RWzJ
/0ui72nbOIYZeAdoftow2My2M8Ls5l2xU+PdeDVrIuOXznqwa55ObU9GMGEuX3Jv7kNCb0c/s700
iaLwVsFRk0nyjNTDQFNWCM2kWNMK+g9EP79naGHJPopN4qwPKBkZv4jfurmz+2/Dr6QwNQpLdUa+
QZzXGEsaRW5TyGOewMYaksP1j5BuKooFmNlAd8XViX5Xfh+RSIrz4UQ+FJI0TkPLUaHhezVsJeQn
T4TfQ0hERtkhoY8g6LJdvyXn1nVg8C3q5S40AV4CY4PKte4ybISy6dedwOO1I0RDHhe2b45JBm54
hNQ9+aAflpmFu40h2BGf+yVxQuV2o+nB9+LJ8wi5lNVpFN9p7aYLAGlNhagP8DcBzcTYL42VgMJS
7Ab9hDUwLqUjRaXlAGlnmNL6Xt+B7qDIi2QgK+tnD9fWuJVrOdknZXOxgFEjycBAGUEdxjT+K4Gh
/viw4ble7+fTavYV0nrHzfrUfwnuA4M+vMShzY2uf+aAkdYzBEh3vSN3D2yY8+C7alzpGtxkjZcS
Yt3ognfLMbRoEyMglH0VrHW6cWzvp/9KNxfp73Vanr9N5ji+P/wb6v3AS7JBC1lIV3FfQ2Pm/mM4
anNEEJpJDRsH39bOxi/XZ58Z7txEbDp2pEpYKVG5Hi5VZIWduVA184uXwJcOiC7v6AUaY4o+uTkJ
TrXXq3Vt0TLCYAHKWmp4lpwxxSTd5r0DkqI3TasjmsfN4juYV+ZnpDEsdkcFUnPi3CyDPxl+2M2D
hicZUJLkEz2TywwiWT45cCCTZSr1Ako26aDvThyrpgiEfeOFIA5aUayfsaHIURrVm2bWsEcaw0oq
kN1vH5jAnuivwqPlMLbBHrdMpZv5d0uher1AKU4jka9fPsyQteunWDZE3B2f+NDsosm542ku4rZw
HwRAEljUidRRdCoOAOYQPllxnSk15S9+xqWXOrrdz6djot2O81U2ciO7OtW7gDIA+fHiIliXNpAv
mve1h1hA5ygFZgW3yeBauyAxUNG7HBcuRw8GPNru2o6S7TjIxRqGLhWsrtrUI4us81LpRz0c+5YD
Wriuva1OCOaEnNvTS07ROYp59prO8SE/Jeq6Ubeb1tahytGkx7rG8cimbErTViTaEtBY6Qh1pakH
ihBWJ5Tm+j98ocllIvDyUMw3gshGIpis0fsyYXU5RCpTG2znSpt5COQHjNeKYwo8WQxYDRUz7SOh
xTQCN2sC6jtDEPczRHlQWigTPShpeV4uoi8sdRJXt5M0PDCwRo1MGBbYhsA3xvfrHhxbTTz0C2G6
jpjyaFDxQJ5pbAjqvqraohK7qcF+KxW3ILLpHdSsg8VvnwquJZfP8NL7vaFk3Deh9OVE3/TmtJEX
Xl1z4AMRM6syFP1X+ONwHHt7c/VBB3OkvW64cTyP8wpE7uCKm/sRg1Fo0/RjW3Hd4n3csKb19jDC
LfKVaY39hwoLmEIBTJJ79Tk7Hq6whdEx056qKWZUuDZCMfICFVfMLonzX0A8gp99qwbxAcYBA3nM
N8O1ajKBjn0z0Pr5L4OaPWJVoK6y9aPRWoUE4e2XdNI8IqB538QNy3JamqJqNAHXyPji7yOQQO+s
922G9isXtaFN2T5BLz/6b8RmfIu8bV1Bk2WccozWKasCbX/8LDL0bAE4wI3xj2FggsIxsphDbUyV
DzUXDAP/8+q8Ecg+ZLgKx4aFnd/zJRSUbNXkpnMhUHF7hEUtSeN4Kf/OzwZ/Y11OLVdzBjj9EBn0
b7IxhjxB1t0GXhO3zwag8UbsInMYb8Ywg5pS50RXvXGl8ZO/NaSNEN7bufnhL+Cqo0EXwvwGZ/6f
FJY5pr2DZxkuZAnN6bHs3KuP5uqQAgz2NxJG97T/b0XN1P4rJXr2+Ufsp3hTcQ3ceyzVyi1ajOnD
FBbuk4GzNV7q/qKdF5+Xyn8k4DydsZ0nHLSwCq5gQkEZwi/ZR2JYFD3kkPrQMKpipH15tK/5oPUC
/GqBNB9JlNzHIVsrvdh+BQH7M76VI4JcWm+hP/ohgfoiUPjNCi1GD41u4G15imymSEKKcjgU6kez
JnX2RXij4ZTZwdQnUQChpVVrrUJ+n68KHLBSIdtmhI5i48vTmvgckIXdqVebpmOHc7hCgn9ffFNj
RWmD7mXkarKfB3+qktIH6kesPzRkj1YAtD4J5R++CjsNJbYbgr2DX6Y6JET/msrVeenasC5fRFEg
uwafsC2fnl6a7AWJmHCsaPvDyYh/lJzGm/Jpf1hA/eSMbxPDw+kILgr/cm7HsPj0gzHlYmYNc2CL
oAKm1bdPiD7qN2QCXwid0AMXNykb10ImmyoSLi17lBeIJH4+mmAQKJ7vS9hn1h7bfycdronMt9a6
KoYeXOQripOBFVDF/4PmnfdfFw3WeKr0SASVKRBB3Yh+uSaai8MfNeBINHH+kYMKL8BhUC63JGWI
V0+O47ttXaiIrJIRvWdyr9OkuiOqxB0TsvkgPIrIk5dsUb9N2O0NCTTKNaJk60/y+Yhu82b0PGFz
Nh64vWtPp+02+Qae11OedZX0TKDZNM0hesDSJlY7Z7Uk5lOKOUiQ8gv/dak/Wks1Lm7auzAzNHB8
plrcj4mEu5evE8kKTFfeJMPmbPtOwIfvgShf9Xjv/LoyMU/IMFnatL55qZA13OavoFJM4jVOOZnO
jJuhovMykSUdmHV6GI74YciFOAQ9SCF7vyfArctelwtHBnNHhXVnvVY1P0Ipj0tEfHVbCBbwuqZd
SqUrI4Im5HibYHmWthqQEdEAo4FJ6ybS68hgHJSgl8Z54NQGyWd3IJh7jJ2wQNuESz3xK++limgD
VMrfD1UTBlSUFWpKD7vs3YKSbBa5qeCTg0CIJyfmhniO5VRCOBKOETfUEXxemvFN0N+xbAcYLYv6
0Pi7hGGJDqm7q2YKj7lw6bJFQehg2OyFhMv5tVzqNS6mHUqsOCZUsKr236/8GrCEcC79MPLdsNpK
D2MnKiu9u8VuqXR7WMfHdkLNxEVDPGLD7Ahr+n/nGzOd9XrIOPtcaXJ1K0zmgkizATkIA6E105cK
83dgL8cas0/D8Q7/Uyq0qFDQaXh7ZjiqEWw0mY17ZV5XJi8QZitfhwYivnFoQkMLt8yj0nr7ma3b
PxHonRm8tGVk0pur7coswyZfAprC2W7/Z1sU5+TYvt2X9vwA1L/hbq44u79yuCJxitUDIkCF7LLD
hDZG/21wVwe7lKB1HGgkTbEAdVQzfJLYlhUSk69U/yFRCbV4TbaryYwWfcEpwbibH8O6DixZwAM0
34uD993Tb/3sSSQWj2C9MugTuA800RcPpC56tH4w/BIFkqZburBVny/4sGMyxNIedWkSLLylV1AD
7FUaeaHihNEzLrtYk+n/QfgTNc28ebyn7hJaaE2jgkWOyOZjO3kNSnfIkKKCz68arUpMv9iOiNb2
ZcjBeCHGG/XGqhlNsEnlVcSoWcmEBxRs0xjhjEjMR0HGiXyhq3M2kWBxbc4/yNKpJ/A8r3Ct3bqH
FbrQuvInehF09SxMa1AeINt/egQY/6gmqXbtNvxgrajTNdZKqUaKIQOUok0g3Ppybb3kz/HJAAlj
5vcYzcF92lecD/LwGstlUK2rr0TadIFCNAgD/c0SYP/IFsSHpPj8NuEkffdofm1in1q9K4zLG4zQ
e+2s2RY1L5WNao+60JQQBcpCy5g9+J0xnDn6EntIqyjHtV9GEWJvSnkY/FLzSA+o8mQXYsk/KMKm
9MbdlTcHEJq38BdXXyU5CTVqpZS0Zosv7zawzN0pGj61+Twuj2LBJHk1vc+Di6BzA5FgWv4v6TZo
XxEOHRDoXVRx3xL7jvs/cXMWNXCwUjC1KkAjV3fInl3vi/MvdqpLLIGZd/s2Lw97IEQud9eE51+4
h85qu0x8OpTeXwAD4f8RpN5Z0GpSTZPGKSUilI3DV+rWxnpJj/gfq3fkpF1UjhxbYqDtqAitv5Yl
PQ6YmElkkp2AzNYil7G2CPXrCXV5K4DNjHP+1nrqJLiMKiqYPsXUBnnZR/z3dumJktJwCIJyyj+U
ltpPW6NdHNzVd3vZkMPEi9W9aEsnvpmNi3ZtHNn1GfHM6mepq+XUzS4QqKEkll9vn8zY8FClrNOG
OB1sL/4UWid4Osbth+gK8qv7sR6jigGjQOssqXqJU2rUeqndxb0wW8zTL+ijHM8Onyzs3STbUN74
58+MqJ1h/ja7mX+EqcdG8UeKFdLfk4YLn5/09N9OHZdpb3yj2Jt6hcUB73xmjKs9I4LClMK7ygzT
qLyGDgprk3+vfrdTVefXHUj1wz7Qkk8XKSUK6R+Sh9ETqNK/52Pb2P2oYRuWqDp3gGkHs8chiB5m
4P35gO9q0z5J3saiYd5gxD7oMU4zsxwlyTF+9xJV/TpCHeYv8cWgqbDMosnd8JRkPLlLbxgLSQBa
7F3UpLv4u3IRH4q+yBuBmkQgDmi4F9HoISFnZMHqfEHRvtRXfBozd17QOS0IxVwqujYdqvH+ZcWX
ULatHVbAIVUfHlqWedYYJ5aSHeykGe3v8ywItcBp75+/x3PNbFqXLq3PDPJQ2rkzOM8xsMgCJEix
N+s/dMupIZ2lmB+Yfyop0GTSudskYWLJ4uSPTmuuZTYUPnkTk4zr9K2aDqfEB1xiHrYdOcMnrldi
0WF7uUrdqK2xTL/e2Tt3W7xcAEdTUkDO8a7Ac/7nDv/LUpGggzzPDp5cJQHwYsIyltiPrcKuOP2X
UxQqcqPtBU4+44SaZN+ka32G5Ys4rP8HqhkacGHqgd3I4KhFShh1mf77az1AiLeaMTy5an4SSoFk
zkDai+hunsBhv7ISbx0Zu4BLAzVEF44ZDN25uM0VdQzbnf1qsdBPKfTrH7fY0dyYsjPsy6xCV9mM
FfpJ5jsQ8hDSolfxTOkq5UOMUIUziPHSs2o6eRfmFlHJ+8OoUEYodhxLDQzQuuZFRzPcYA1vvLo/
qEBPjB3TE7pr3WRatFu96JPTIZbviQvbQjttK2tHAgEeLHdOI6htXwesnYf3Rl5Xr+sWzi2x/ogN
+NPDbvbPmllmMf+zTySbtaE95vTnH4nkGXik+v812mfiNJKzgC8/QNZd1sAle6cniwOJXKCY5BtI
gn2iGJpF1VO4VeY5XY/yRRyer9/7IKWOBawmvGZJNpf1qbNdrDMuflfLpR+6hIYgGvcH4u2C6tW/
hX7qNlVgqSrnRxZux/r50rjrUa0xe17OWzpOHlLTTaAfyilo/LTjMCqWQNjfJtJnqlH8c5EKHB9p
EjbMmmqUZJ7W2z5vubaLpmpBBq1VMOjI1OPPXOXEmVNmL/cxxArMYpARHFvP4ZU1XOHdWH0inyY6
BcJF1o+g1T3O+lcZEYcVN4vFRz/8ahi4OWNcLJEUSKgoyQSqkrsI9CY5itChpK7SU6f6YgW7Tq2w
V5m/bBtD+yxr3sgUwk6S6KSeZkcMmDkIQ9V4GuVU1R3jFO1bVLBMnST8CpwkhL3hMnM3mQx9SLz/
Qrkvz2FdDXLpoPfT0YnH40xLRodE/+YSnvFFuBGjXlsz11E6qnki+aQaJZL11fA2abbo3NR9lO9H
YsURZuH0e80m8semLbDD11XJSh7ySdoXWolpmZP1uEPvfG1sO12ItcCrz46Qa7rQCMIk/o45mZHz
mTJOQu3JXjfn8jQQmGkSpEa0cRw8epNsDbYNTugWZmvpwAcDJorY1cNP/KrJQJI2CufKTWp1pyF6
XZqo6JmWYD7UrZNfXvferNqJ7aSFwTr2juTPPSqvepJP24aShRyLoNbx5ON2LEVNfSEyii1TNgkd
AaO0kCpP64Ri3TweuEtEe21pyjMsBdUrNesQ3VaLIZATEqeiu57mnl1HSvkzmtCWuheGPWJ1V29A
fDLLTCOv1x4irZEd4d6vbmqz56yxngXP1ymbfopdKYEaAon5XHRjBiHJKiCXoXSUuiNbsYBlA/ua
1hO32jEhvYsRB509uTw+oDVY+lTpf6fMOns9EcmcHElo9nSDVqpWG0iGgeIQwsR8iPxMhM4PgWeo
D8LzF6dMdRs/xGKHgE0hYtr5KowrihzBPhm3je57QoWF2N5pUDDcU2cRfBPU/M7RnDoZU0O0lDeh
4Uv7ElTOtX2nERBcrU/vxuFQZEQOGEHjirP2mXgLBBuYi/30hAzqLwfnrdcw2wjYsIKBymIGX11H
4DNr0eQQ9OsMb3S8PquWZ73p3I9NPH256z5WdNXQc8ukTk8ipKt1icfpXL3GNdIAKJohFdASIARp
jFS4NqtbKolf+S6senGrLHAjMHpRquncWZ+u8Shoxm0/3nCJEGaQe9dSNIU+4424mrSDoAzS1wyQ
K5gFt4nF6b+To5BqcWuEyWPcCcTVMp/9auTnOH7635sD/bZpj0JsyfvYtlDgfQZeCRTpxBR9pkuR
GySyOee+iiOyAJHwS1douXZp7PbGysrifn/yS9RzwhehkZzWUEZVErJ29NkLOevQs7qOSa2UL1Iw
NmeI/CGL4pUJxXeobDGkAka7CNOzv+vQM0C/7UJtNO9oD0RHaPdRsVY7XZc9unZseg6FFNtKtwTg
McNPBn1hNe2CPnKE7UqOIwnHD9jMVXJRGTV/jLnm9qvUc/B3IrxRwRVtXrTZs5kVbUTE99Puqn1a
aC2LvxUFH2uuX6DTF0M87/1Chbt+uzjLa0fVoVtNlKgY+VXU9XE0nMEkKpZRfUsrxJkM+ZwqwXEd
eao1ioaQ63/aIRHDoVo4iytofqq+Vf30lw1oV0pTmZLe770LcIqhaGErQt8UVdES1pSMs6o8qXGK
9FN5w2vT1PMAffeS6MFiEo16a22+yjANKgHXQnVRBZCq/hzb+l2MsPocOV+93b75ePKBwDdMJs2X
CN/EfzkgZROrfjglAbYof9Ly5FRLDf9OKkskcYCuqB1QmL6FWjVvxWWrqcg1Lq61vTRySZD8CsKM
9tg0C0TvFUt2JBkeiknX/ZvClS6l4MP6m8g+W9t1HxhrGYisywR1jewslPeeybSNJVvFuj3XMMhB
YQ3I4bHeXjq82C54BRPt91nNFwRMRZySlaqq9RG32MPEYhYeD84273Q+S3tC2WSlF+kVrIV5o5JV
9byxWny793ezeNl0GlwPVbHQq70SRlTHyXe8ZX82rH4MDKdtBxZ8jQBnuxf2r2nkfwr1wbzmjIdt
UbDw6/ObtSL7uN1kT3rTNlSHfPvLRn2+3pn6gbm+N+iM//vIQto0yPHrLJMrnsokpR/CyV/zXlsI
MssfhzRrrN0aZtD+pDehl9d2W9iBkVd6SjlegSX2/rF6uNsLHEO/686kRuVC99QOXPiHayP+5D/q
QWABn3i+Pzu+zl/p1D5hWH3x74xoc+VTAWll/ZeYM0d4/lDjfmKTtyACIddn4L4xjg992sEetvZ2
ebUm1Oc7lY1cOyh5J3yh7/cSvM9HCaH7sjtmRMsz/Ao6K2nQYxV7FzcnWRr96HncxnQQ0ajf6O5b
Ej8YbGFAwQnXFjBpQr5L0I9/mJoNxS27u0LgA4oKRgzHJJWeyKBJO58+nYtpyd+P7fCBOs5emJNM
MT9zL3s+3m1sDqLevXUusL/O5Knvc7f2IxAb2WfAeEg/HH5dL9/Y7JmT+DZVKdM05c9UJGuEGHn/
IcyKV1muDRomXMlxHLPf3wCdpLuyi6ke2CbVGwZvsVuZm+pPcleIA1uGTvUQ7jBhVdswZIelkAiC
5FJeUrRVvdbNBPLdPjhEpaNb0PO1+K5PjttTK4EKnSS31i5JKPrBO3iIK4KJdMlBq015DdG7NpxG
rqgkZwbMcOK0NK3j+x27g0sRMMYDib0/lpd20xsxbkEXs7KhirV0gskNDtgFIHqODFPREq+JQrIe
fhGfLV/Ru7sK23zAl3/h+PxEZSbA/AbSbq8kRyjoXdiThRCZjGUG997q41tASY+4GemrxrdZUKrZ
0IkxhdcnJ6MS1h3cINU8mqOwhD+jOqU/zksN+QVu64AMPJ4bvWx+00zHlnm8WNiOHFNxEde0Ersh
L9TWD9F1gE7gwr6skrN2Dj7MJx7cbNE8wN7oYbwIaunjnzJOw5XmcjciBqbcVRy81EAQh5sg/Scb
/1xg1wHLW0au1hVOmvOIu7LVwgUoNI15pOkwqknZPOL/hnVEvUvG3rbtjwmw4nk3foP1OsVRcIxz
7u5yGDMpaIamIGdQs0LhVktC+ZoBsOBMj+k2ll3/uo5PJJ7KUvvBIDcrmq7sXzAn1Hblc2unHpjR
fqZSyHTLE8C+AIfyvSAvaz/4kS1ys8ba5RSRy0NnloKNpJpZMrG5MWhEgGl9zjerDYGERaUR48oS
N497zpTbnWhY3loHcUr50wMf5UH60FMFEnlbov9eyvwVjGvor2A6hPvlkKbI5okdtYHNzM4QfQ6H
MIF3T50yuW+9WJ1ETHsmmEPE0S8UYgZ3b8TR4VNQyeh26lKK9PCWlQcliB2as9yhGq6fX8b1HcrR
W/IeuJbmP5sVGYWAR8GkQOosC1tO5Wg3sc2yaXzYwPjnIsu5oxMb8YpLxwJfiRu9Rg0PBdzTysjr
Zx3fpMxWFODJDVPYsnR7UvdVAhsv0ZFEIyfKQEjO3h0EQ6vdGJSXeCoGU1+jMZ+A31z11go5Qr4V
TuczbENzLdA0jXFxd2b9gPqG/s7rSymLlXF2PiCANMaFLdUWzvlUZJitW2/T5CLgVRrWwxe3/XJn
Nk5JzgKTna6CLfBnVjj8i3BAHH9U4hXV2FAVRh8G6ghf2qsUpuwk8sXhp7grf2UoqUezWAQG8uKd
9SwUK1kY8erymfhqDLC037NBxCUqZJZM5MTkXBkZjLGJg0AwP6jyUujCAZnwMT1f3Ng+JalCFGj9
pwThE3wHZo85e6e9fpVtuINFFX1Uq0JKZo0QmEOLcsIGybgXSTe7llcoPd5aoIQ1QkQ4rwiafBH4
Niu5qsFjwK7EE73IYuZqK6l+kK4LMj6HAeKs7SSBwHUQ6Sk+BiSn5eCC8ESAdTk7rI5ceKDSRUpC
VJ52RvkFII2Ioj+GcdSMqBHG4QVE4lW3E5xkRh7Pm9reCN5UzKe2bjmEiY4oT+MQn37wh6nf3pOW
VWlzsxgvXDRC9Xt7YoLoYjqTyXrWHPgqM6QAlXQBeNDQzoJiZjgeUpSsJQbFImQxw79dJDQ3gLu4
7GkVczTjUvjxmmchuhXj8rxw92mP7+xE8nQ4yplaB4ViUkiWT0GWp0gYQeONOQM+3PrjsuJcTg5V
ZZT6AMiVOW1Ge1jvskRpNA4bOjuBEVbO58jxoN5aAxORvK98uJHekUc7yKzlvTJejnsmIGx6lb6B
dg6srGQm/JXRJxv56rpiCgsFz3azC1hlyb2ndE4Yp12SQ6EbuEVaC1LkRQvaEjR2LawVRARRt8sm
EnTXqQwbbHUEMgrhAQUc/s0rZqGjahdS4HDdzfc0+YIMcByViQqzSw/Hb+4Sabo1FQRneWcvCa90
45AmOSyQlFMOpzl+6JmzYAx4MRFcUz87TFXgvBAnazjGkxysqD8HqcLi+BfbF0ahg/6/+V/4V9uo
I/PCW6eKz2DikRI8WQQEln2Uz+S5Xns1zHWBAfYMF07tj7hR0/VgTPx8s6d7zV1OO3TQoLeG3UVl
AjlNaQxWB4ZML86f4e3uzK9/Dr8snigCV0MCmfbTC/6Yn55DKIo1BxgfkmZZGsCPKAcNZ/rtxDCS
GQazDLpkI9n7HuXM1MsQcwprL0CG4KwOyfo3ntDr6NIsH5wAy+FhmES4Zrk7d8bQB44VoG/VkZa3
nZZXun3H87PxnCRxr+8NnjwDdMj6sOu/stVe7ycXFxtQdn6KQ5y/zAp1rsAVIj5lpiYdWlF/JvHO
Wb+tk0uKrU86efDfLt3psBxFVhVgZAzhGkZrj8gU4dPnExGaKV5Fj3+shwO/cSbXa05t7uWWaYTL
u2U4eEuN1hDAw8jNIGKYmBAFITBwnaJ05sKdSAZWZriHtZ4e0xUcJjuIEl8u+rg4miastSnFZaX9
MRGZqN+eE6asqjuso2sg5A70maK1iSru/w3a9zLmjak69Vuh6W8zI1SvGoyR3H5oQYsXaaGeTD8O
5Vu9mLExheTPYWioe3u9kPv6+bjFfWgytHHD8UeA24eTwDOh1cdJd/xnYKXkgbT5FNJWskKXr1Gq
W0x6DFoxmtEV9jInI7RHauyzNngJT/BeVBOu04EoyU5Q75ilbP8bBbD5rfaT9GNZNV0tI974DhtU
VzGIUgw7mS4QNYqkxjCm3fyhQYoc3atHuk5mF2QKrbyfj5CSaL5bTXucQ7ZvEgmJte0cLAOyfQ9N
IvGoP6wapX8kbMJ9kx5RcZ081hCO6WFJ0RzwQdqDlpgVIbnm76KBXO7DamOShvboVwto0oQLkqK7
/and21Np9oYvfhDLWERgEU5E7yrgqCl1eXuX59RLHTksRnpvWKVzSOkMre6TMF9Tc8laeE2KEH7p
Bsq/sNlb9zcVGyUGO/U/k0b6gZes2VMeK0Bj2R7KR+aaGaxDkaeg5IjNXOJkba5oioPTFDAaPDNB
JZHf2jegAS5+1faWPraSvZUU31AlsD+OU8oeP/QvWEcamKmyuOq1Sw8Zf8eFeWsM26x9T3xUV30I
bOGhvRjeKtgf5UaRswpJDtowfcZ+FGGYupo2JcktKzeiMuF0FolSci3izr3S+o6eDyDo6s2B+Ukj
EzjzxQNDeLSdnG2qs1z0zM+nA6ZPaMHXpEVX7Ya7AHdZUizgDy/HNFjTQDa5DgY9IcNWYMGaKAmd
lfrkCrYf1jnsbkrWRcfhwEKuRgT4JK5TFbfcTDGsB4salk2MWCMtqmzptR56xk7DBho50meyknaL
jbde774iBP44UaCrk4nGyHC0yhDh3nqLYuTUsc5sV7sYc/9YvKKPYvS6laVcH6jHLVdZBhZiWlsf
B8vmvljr0RjDVTE+iJnqjA7WOq43ikuU5rw2C6/HKUL+DvqxqJdI4KYv/NsGhN+/DBwWSWriQz11
N2nWTjGPQySCoDSJtKlxJbrP0E4DOKPWR/CxA3VaElARgKxUcGTo6MpCEkfTxKg16RYZIORIhTMc
3Ay9C8FQU0zNbiO76yJOmK/nHtSVgyW874rjsiJLKNM0skTk2aIhPK5KSdqVGWAfwzOboUnZmiz0
A+0Z8zMZ4tgbKUTZX0QwZGEynTt9wnPZMfSOmJxJOQAzJYfKJ9IIZS7aynDhL8U601DeMKNuWxNp
sIXwgbZIsNRQaaStiQwT6zzHirp9DdGb+r3JvBP8bBQDgErK650lHk6AuV+tXleT8ojhgWuYyvNK
jnoHz/Wp1/nDzCDJDLNNb/vZyBk4/PeAolAUmFaF2gOy07ZaP+KviFm1nKFK9+MYKgbifcWP3Tsi
EVNNc5jmLd0i3yGnAZrsfKgzr5PxDsPRIg3DLGYq0ojZQD9pR6szugt2JGnXhrUjAtvhDTtZikEs
mxXe9wEBqT2x8xnZ4PSWfS2hl49Ux4doHrEcvWjnxEAV4Y5muvAcvO6bPBzsF5UuLTwNa3NoVbHI
UfuvzE8n3iCq4sYjHyfgGQBzAOIrWISCUr4THCx180TpkrWkaNPUkcq/K/afaSLdAoEeCIeF29c9
dXxdj6JK+7S4/zLQDOgKhvTooJGmp3fJDR8hyG8D6E+btOPqymys28P14Oil38pjN5gS48Hinju0
Fc6rEkfC+x8fXpYdvK150UjPRzjHgIHoj6OKWeWufFEt4pSdp5UkMWyzC7hgqw/hEHJ/DvN0hHEJ
u0Y2X/KqGFVCnMLlOnbV6eJ1lWNDM895vHQwE1UqzZKIZ5mwfcJgE2xLlOZXMhjZSfJRnnUeTkbM
48Ekpv4qyS8BBxEH0L3ZQAUUDSlg0/KkDgUhflUTHj4Nh2eElHejEE+99RQUE5QKpBAKApRGzWF+
BNQrubpYdTsx/V32ELE6HggZi9fpEd80xkytUYTbwc6DvNFQ5GGnwbK7478DMMHW+EHwFd1k37R3
Oxku9DSkHat4ld8DbucUNy8dr9NS+ektFxk8bAgXIW5Y0RnsDhjsAs9ZEsjPfBINtilMdn0RfNNk
DkzoHQ1z7jEF8qai2VvYkCIg59LEnYwVU/AwvErrrI0P/ENkCZtlmSoor4dG05lZTyaQPDBBKUJe
20niPBwh3GNDXPCvxMNLTIFPVJjgVHQbGIsL98BKFREQIQ9RzDfPF62F84WrF1/D4UNnUklqgbjx
UQhFVe0B0aV0OoRNeRkJgRtxCgr6u/ITNOAx7mxKPziWzf4dLIw1LTMHLPk1KRTMhovPY/rTXmb+
gm/b+aVLBrLFbn6wZVW4h0LV6Pfpn69YcCqHPN9w9FIjszYO15mvrI05L2KQCfDbloxXo4ASGV6d
0G7bmS0ksywAyOOMO9LRkqvcaSNrnX3gihkjBWL5/rCa8sNaXq4Z97R2zNwjRB4HMreiEQgupoPE
wBgThcpB3BZlnx8q0KxiVEWkbBgA9Lilbh6J0RbR6eh9R8PshFt8xoyV0L8jQ3oRT5FxqXP/Yz+Z
uWtuOZsovDtT23XzqPT3Ei5SgU872LXUudmzvslWFoIHUPxJIKM0QO3l0AEjqdxAALLClVdBAEqG
yHkJsya7OiWrThH1l7tt9ZXwdK+EikvZKwBvVfUkqSafLk2QqhbrWzgKKGkbwDvU7BezAmVKq4b4
W+2vTJXcWiG4jSwI4A6Qdx2oo+XKZBkMKKgoBvRiIsfUVajOE5xNM/3CGEbs+1vRVg+Tj5PbaZLK
i0dOqTRZV3wI/TD4U5NqxUPcWxLa6gt+PA16m2UmcxOOAljKZjHlzCkc2Fus6IoYtfGsfeOfm5wb
rhxw+h08PbYkxh3kLXy1rPOKagp9qLKqAGUB6fI44lnaREO2xwM8/soPUKdNxIug6MQ4cTkOgO1Z
up5V5HedgNFbZmyxKgxQc4jRfq4L6Rfjot34PnGHMI7IXWRaSheX8Lrq+2Idda1XGZxvvrlnvAsU
exLa7EdUmp+Ycsr72SnNbMtwKTI09l31yLu07n3cHp7x5g29CnSQIiOfuMvNyovrmP0GOqi/9WMp
n43PMwhF+HY9UksPNma275LpmGuysQ/Cg8SYIwIRzZKu2Vkn1GXh5wvpsCZAQldyC5QjPNefy4j1
YEkWjGgGw3pMMbc0SlmUoDtF2AKiZfexXLJZqOy44TLvDVMChiMTc78e8isLPhZBjKx84qO8dZlt
f9BWhEeqqs6cu2zBZugF/xX1E2n+KLfj7Mi+1b1vwPa9dVCuC5oj5NcDV07WpWq+Y06bIzu+YGd5
VI/7S6woAPcncAH1NdtrdJ6rLuh+/4fOMkSOmrmAmVLScXfwIUptv0+EvQsz0a5FAcy37acnB81x
/JL1HtlodkTmmbIvaHlPpGjUH20VWZOLl5tKTI/bp8cuh3eO1nXzQFh3VzULt+hCkTYg28lwpDcg
4gjQUls2eZzUUBOyOcAN27Ws4ginZTE+VM8sAaxWkIDUjdnmrYnDC2ZiLgavdbkIkytkJJPQiPf4
ujORw/SaWHebv1B+L2o97zXPLPosRDvuzxU5JVDSUeNgLiNPerCS9LyQlLifYEA9i4BsNUI/4x00
96uO5dK/lB7kbEoZcQU2Q6HtaLh4jummY07zeHzU2haN/mx9RRW++aRmoSVvViVROR2EAo4JcZLQ
D+IDrGXQeuKKSnvzWJdWdOBujxX6y0JzWd2O+pAXcIMyue2KFiH1QbPr9bwE+KY7Gnd56DVcnawx
1tnIScYxbEUmfzPzZjYKuM1ypX7p8o5K0E9BxI3KNEZLrvijUrOXXrRfHTQCRxf0tBYwajW6TCQK
W1+6IKi9mykDblPDg1CL6um3HvMM+mAPJpnh9qtXrec2kDkjjocwxClNhWAmHSumr4Gs259zgKWu
1Pgy8SQV2kKy7cdR8wDM1fVHKulgkvzZpxdFe4bYG2oW6xAR/ExAfnEdI9t3kw3qsKEjx65iyOBj
zrQKtaTmNwnNmWTgGKG52Xxy7CY8ndfuezvYiX51go9415qEF8eG8fbwnrryi8y7j6EVm5EF1Txh
D23btZLO9Cdlp+otvaZAITHXZpsWNAw1QRIBpnX8rioLuVr5PW6JE9a9iSkpCRB3qB9rF9UqcWKE
IW9twdsxp1Bz/3ghdS76vXf+aYLzPddU5Uhv5zVqcQoJKIdTPvDwG6qus27Z119COb7YHshNReU3
IAzPXSKQSxP0jl3Tey7z+AB8+NFe4gsXKaH6L5tEAu1XtT00iolyTT7+TwyEEGo9gf3nmvQ1hLk1
lSdk207KogwcRVTHCN7g02wX3enSNu6iwLOs8lf4+dSiSuhdK9az9bGgty1O+WF/M7kNs2hvv8jl
BXFz/PwpCxlSfB/j/2G0zuFdwc31yZGAjayiJTeqm7WSW3PkXiGcgD+IOQJsjZKAcVh80Ggg1E1F
nq3kE8Yv5kACWx0nGiMowThoPqZdVhLX+Hwp7OhCMopzydAEygiJQKQOTDeatu6RXExD0tvAVNHY
w2cLz5/bbpHlub0Pb21cZCPNx44hoEJIZ59k0WDLsR3HJhb8El8TwiWErc5qAcSkVGXW1tb6kuux
NvCzRcP/yb9H6FmMZKGmNC2HeMMNhnErGs+zM8yTQ73QvEJnBgzb1m1JzOXnJ8QZOK6PrSlPB6Pp
JCj2t9qkGSbJ4rlS0vbJqOsdSVEm6fJP+xECf4DuVz6s74hQQ+AbCuvhJK9SgxAKHSwVdo4vEebe
jrnmWQrsRoypM4Sq3BMUecyJxDqa2/UrIJzLS/GU9zMgzkfLl7jyY/v+dh14AFsSihU8LQyfw5lo
Yod7bPzfp2pSVmiY4lgGBae/iDNSHo5LyrgTofM+LX2C8hn4/H4gGRuJPYIBywrCwAWdtrJ3Ndul
hgSoNwMY/ljYEYUJKzM1A1r+ES87jF3OHBEXbuF5y4V2yV0CEu1GgOW1O2chGxHJZPog6L4B3a1E
BBrFLaoRnQf0c233IYoPeY8gFCb+C3o/005i2KIUo+NiOZ/JS8XaK9hLm80Q1lwdvGXhwy3D6gaR
L3xO92BdkDg0JisRUm8cojxuOejClJUrRXPvnd3gmetidCPePGw/hTYmyiFRY2hkAOlrqZljxY0g
5B+T2SsM4ryRwTV7tFgOXjgfe5ibaKB3xRq9Qr3TXFSkQx5pg2/w2Y1Fw28OzYK9zGqoNVPvzHLt
nvCyw+h3IJMNJq4utwuhoU5H8BGAgE/iLPYzck2yiXxYaV0LP9Qd5M5wjJ67s1GI73iKZGfkoBWW
gUljBId1Ea4jrovHrXerRNk9VGmIImHiuuyFF1kU4R2trHEKJFnE/QxCfhZJlNyHReScyC5ZufJk
ZHbpXDztk5TeDhKA/mlw796Yrgsnbz6bss/22zbHGmuXdow6ZTdyC16uNA6mUMgDU1U/ygajk2dr
sJY4d5LOrI4hUfT5B1naUFzDNruHmX9AhB2/HpOjYBzNqrCSSeJvb9WtBRBxtL+6TofQb7b5ft+F
WqPrGa+tsEOqttuYYSTTmCtv30p9cQ4HXZWYlVU9vWnRd5y9lm0yCN7eRFumjSPvO0KZqvkG+mbn
i9hB3Q6oqaizWY9cW+LXM38Y+o+WtJCzjCK5lINzQirSmaBOJJilXKwAzeMTLN7+Wj9CKXTHXpa3
ic/ZBld/lO6hQOTvNeAfse1UpnUL+IPB2hKQ97MzzfpSpOr//Ukj5rq4q8hiHTMcSztxXDh6HoF7
K9O8gPsfq7qn2osumoxy4KVSw23OfEoT7lpaPjPEwZTwtjpy7Nj/XtRO8gaFufHx1f01JfCVZJLs
G8FfnB3qLHLdqqu7O6ZrBbN9He0fAnZ+2DJDH7IsbqxmB87V75czgCV5QsCO6i7Jvrx/W9mHRXcK
l+ZI0zUsxza7GAGQbEP0e2piOjumcaCZVZrMgQb/1ouhYF012hQxX3UpGnM3uwJ76oKT7DZcMmXS
Abnz1c7mZw03BIIlPsPW4QY76NagpNFrbYCs/1b8FmY33UzQ2q0AZIlGV0TgCq/FDk/Tyr5H+Hxq
j3xr1XPzz7NzV9FTdGLiT2cI9oTsUeZFhqR7neg6ezfA1kvriuLFlr+DSKjyoVuq6jRccWzS2rTK
+2ZgCkfE3jJDswkx3VePhoUvZwdRv6rBHkZ6bT9oGEGrWjbO8fYcuRGaWa15Mf5dp/FRco+JMO/N
nRUzVQ6UXcFiHbvUlKNALZO6AZgzutFpvZNUx9xrgOSpTBg89f5t9/Befjv6tqXD5x0UcawiO4dW
sdmbqdrDXOGPW3IyXMJ/SNaYGQ+z6J/qPnJr6WES5uFxK38FtBRSNnwvZm4+9ClZ
xoklfmrLwfc=
`protect end_protected
