`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
G4wGkNrS+AIhYE79d/QTzP6NhGjKFHqftl6tBbWx2crnKKUG5/cDUSxnaFlMm1FzzyslqFsNa4A7
YZFiKnk0UA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mA73bcipAdjBbvSOQ/4ydGnIKw/PTl03myG+B4a1ylGfXmpLEyXq28ZrYIT4+GulBFaothXC2B+f
xAyZeQiq7RFbkC9o5zFyTdRop3r+Px/dmg/ly+JXgvZ1Yo3ta6PX8SiMAn0fRdCq+OCLhRzUPytU
fvLhPxg9OGY7E46tGiM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JOepBOpaP8qhKb4hsBLey3NK3kRm/fBLptS9TXya5NYt54bnkYGoG1of+GULev/0H6ncoVN5nSUB
Vv5lGgAJzdFTyoiR6pCUULsmVisojwLvua3GnpToVVCcgXaeMZe+OL9YQcdTh1vj2dAWPNeskJQ0
lUXQl/KJi0ZNybXTFvSeqVf5Mi2ZVZnduD4MwYlsw7rnzAQV8ut0nntGhGcMkDXCoKoDvk5nCQMn
U1Oh2O+JfSAFYHr1wkljRYtF0Af2qYfZI3R2YOZzVkrJku9JzOs28x9W3kv1yMeZPfKFoa3fC8zF
ZGqALqvyQLJ8bP475TjS11eslPHyyRyUz+BfOw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fRGNdQUGhscpGarB7NVvvnNBMQTxvOQFSNMkBYokubfgNfKrRNytoF3ilxWsRp8vKNlfhHjOfztX
8Buvwl7S4m9++1ZCTp2Wk520pBVZYwC/QMA8W1vNlx1SHxU91jxt4TM7B8IDS1XjSeuiwYwUg3y2
kTeeftPXHeOHhWLhTKY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CgID+rl7/s8nf1Il1nsOcxK7DuoS70z6QR/xLTpE1XNZleurWvvkP/7mng2cmUUpvxGujNZZIaj9
y4QLtRjVizsOQjHPpEbGre2L39cSQXgATPEz0LWFqwGood4XrYJyBv6lLLOg1oB+bi+UH/JsZB0Z
xMeZmRbZZ9OLRCvGc9Ts4uZSjlVkr6kDM79hWheiDyHiOOc9O8GNQ3DhNJ9787YLfHSkYqj0GkaA
pbtVdLq/ffmB0SsjKAjIXY0ui+zdPIE8MRpLUKsMYSwbOMel+uC8fvy7Yq1ukAi1w32pudqdXMA1
yV255T//TWRVgNRyvssaEdoDoVqRvgJIwtWZfQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17568)
`protect data_block
OBQ5OurkCAHuy7RbrvHHrQkaf8UQoCIxWza2maRhwrPWBxbwDEW72RqjI3by+0UofQX0bRCUFYea
YNeMtwBp11klzXNGu8UA1nuinWYqw7FaD6EId5PfvsVkNFZL7fskgHZHTKA1oRC2v4ME7JXV+f9d
/UsF4IzVQfDh78h1bx3fLWRFGHC0iwbnKMCFEvXZiMRrMORG/D1Yv8Qwr1HfYS93Mqvh0UCFC38V
ZT7cIp5Y2aZCxaGuhQqFMzqWiRQVFNhwO5pFBPJLbaH5E5yhDnIMnJdQYjEttUZaYh5cuInAgBAf
mvrDmnl9b+y/FLC5AXdHTEnkIazbcUXEUSU/Hvai2I1Oh9WFHSWLtm/aIQfibMZwRBHKYdkNcS/9
HyrJ24vjWxr0x8hmfY856IlIA9qKxCdU1CMu5u8abey604GErMnka11lGaJLYBoUi2eueDMf5hlR
GZav6dRqdiiEG0sbqo4Rs8FmBf8JZAg55v7sBijkeD2B2DiKDsHFPLuWAo/BbZPgqMAf48PdNXZ6
EGtWokCSw9pSjRbY7JRaFHPe0OhMjjnuBdSxC3R3bzrQ+/E5R52NkN1z2rWlklxXFbyI8y3/wZN0
FonUT9z88CkdMuWZPCuxdW5MibIfl5ApNzqlX9SMJWneE1YGBT12fEoosUnNh0wUUZzfl+BABcIW
KCE47r2KyCaxdjaCzBpJb10Q4pi0htu8BfD+tc7OdIMbxV+vULkguh5h8W6ErG3CA6NGtQCe0cbn
3ILu99It4Xd+jmc8U9mlkHD+XVdC/xJhcS65KS0/sgvd0IkXxcx/s6CNdBN8qbjww8LRopmroF0w
vvbcAmCjj+a3iMWLdtR5IAoZyFP7bSwuO6LsWliEzoWCrgUyJdTl6cjfmIvkFEBXv2oZM2YF8MtR
psYn1MUVdEmMoV5YQAv67M31/hDAcnnUE5e0zqV8teSQP1uY/JxLu3VYrF4/NgmdlixfaVCtOsg6
mU3hitvANsq/wjECejmMtHdpL1iuA6vfR6kv0h5Fa9HF6CQPWRHgfCqoPxJnVo+UsDd3+bmNfAdV
uc6/V6mJIunMM9ukcvxpSxnvNYpThWEFS3hJozTdVgLcdQbIVyTK1YNqPHkzlNA8O2Z9bcFI1ADA
gH4ORSYdHRoKlLkcyXzW4oYM1V/TpJA2Oa11MH9XQtPhp6ldH3wfJtbkOJW+uHuZdivKVJT67/rN
WGj5bfMa4ev1VbbezlPuTlwdfmaDULhtbcPON/D8eQrffDqnhWAvqN5YVAEVceBu+0o6V5gwtW3w
1YpxOPJUigT0HztRGcpBB94TCC2lohQi4ovaJdO5hbNsE2WBCX9/8KpvrYI+EmroRpGeBEjqDwjI
qgO9WA3XsyXePfT7QGFXUFdN7xLj9d3Qv/5Kij2lv6WGdQjyiKZTyKOx2oLmzbAjp7DeoqiYJZ5o
fPsA9bY2j1MPe9mmVk5Wci3BNlhVQYvoP49UMCO/mAx11/BTVgi2YgNepUkD8hlDx+Kr4+JUhtmR
TelUi+WgvulgRHFZNktEckl3EvYw8FZ+PTbcHDSLLVO9ak+a+otXmGUvdArAmGGiWIBXXpktpPIb
E3NqF3hmF+ESIFM37SBYBuEFIaoG33vyUvqO2mX837grh6uMjODE18lGZr+LWDwy7uoWXDE0disx
eIzFPndggCxCIqVpZkvS7s/+vmfK0kV4Xoae4ZVhqJXu8qN0zHBjVgqGImJNCObR7ByzZV1R6OA+
A96zvi6eYZRCraVt3Kx6eDjRY5q5Mo5x0CoKsedrzagn5qHpvBKh7ejCQDBoTys6e1ymaEfLyegH
e3YMUj0FeinzCRgC8b7/mbLUnZx06yg0jEnC9aDCAG0blE5AAdBs1fY6yvxFk4KpE1DiBNvrJKm9
wybatbU9EqpIqPAnwm+EQC0DnJlw8c1MV7m0cR1U4igHoygYNJofjjbgLMloiYrhFsp4pOk8NuzO
mC2nn1OPjoBdlcHrqERwfV9AG+05qerGEustO4k//ujkL1b4J9Dw/2Tz/8f3hzn26qz6Yp6E9fsS
gXWATcMSpMp7dcT51xAYS4zahxbcPs19GGHp9Z+Z7YDqMPzgiux7J1O842H1zlvCy7Uav5QKyUW1
Wz5KjmKRYyRfwV3acFMziN86SRftlb3GYfqa+dvxBEEJMGsDlP7Gs3yuhKZ2R0Vs0aOzmsSfMddw
xTQeE8J745DDTYN8ES69wvcW0oiljCfXyY8mU/Z45y1Vk0TZRe08LCsruXATxDKQ/uWAoacKH0tD
ZXpUlqRuBf/dNfuBRK1BBcrK1EgtxLaqRronZBxBCrvy0GDXIYR/+MjHmjuUZVw72l1R8FxUZb23
jQifjZmAY2KA1BFPTkVF3PTxOsj8ELqBlGFqbq8Pi0MYzRqK/pKRNczdKOu8LOHYqYXAGBRw/RxJ
7082zC0qYsCExUujI8H2o98fDXPH0XunyfxaLDiVBz9HfPLHocewSeUJTChFt7ZiOawPnsbMrSCX
1hxwgV81jF4fY7WHocYoI9HuJ/PPNg+1AhPx2bo4l/ug2SuGlBAkkQaVawDmn7lRSo/vSEM10UTF
c0em2uq7L4dnDNJXfou3x/ORdAi+jmC9nBnNHIWCaEmfO+Hyhw3J47uiIfm+IbxXeAwc/VdVeMTl
Dbqh1eY/BSu79P1ynhr5ru8EWFGorTuOZ8rlx4nnq2z+nDzFE3rOr/I3IEzUyAsCvbpN7aVgNXZD
FCuHzhwtPljhpCFT+ft0fZLDU8kxGdvS4EeHeGx2bQVGmpGRJjNh8x2ZWmcFYDHEvzWaOEjRMhnh
HQ5B4Dzd1IEtrG0DCH8doiux4i7+xhBw967M9jvuyz/Ewfy6UFpWC6pgyieXgiEv1SzVJdjcn4Cp
07Ub/ectNVD83lrDLxuhxlAjDZDd2z8yNvuFeu+2++CenSve1MlFJ1VMv8/5e1OW/OB4tOJUoPy9
iQeMMRxzmcP+a92Lzt1g0lE6+PvD4b5NhH+A7JVruChMwPpFz9fzpV7jsB8tcMt97n0ffoaNtOTI
VQx+/VtYOLQiDi//dGvDJxxCBeSvzkBDRoH04/SdHbA92ccv4RoKfobzpR69W/D8+T7bvu2vFFZY
vpWwPUw8gVPqHmP4TPDTiBAKtHN2XRnxWQZVbk7ZHYDTioMQeZS9scqWsJQxdVJ2BzIl93JXIz3W
thImdtxXhATtFFHXHQTR1BEGVyZWXc6IMyJ2xnESGHw6OjSFcHYDPWaS6cvEBtAtAeOdzkIy3Ovo
FYCQYeEg522yK1vth48XuCGlEft89SuDykxG5eWjPT/xPlFRhRKIrMnlNzu3mGgY0oDaNNxX2VEo
9TCCICzNx9ZKR6A4BMD56zi4mHv4K6WT4Uzq1/oZ4HNaESPVM89s5BDYsh550efATK1cTu8Gpw2X
2aBNuhOcjYeISiW3JZmFkOeWIAcvd2lfSJDIzoWlMY1K5+O/tVJcQTFpGwhOHKF9oqd3BCginB75
j7l1ea6jacQPbUVngV1NenR2BZsGMfsXQPKe9oxn+BkO4DOoxEneVGQd6UF6OldMpDxZBWpiBRy8
SSelzw5/44puI91Jh/VsUHfhFDU0yEXHQljHBegwbJVwyRnl++SMlOlX6HcZ5kLWP3j/yTDb48ev
niSt0rDY0JmoBz6xbI4/jeTkqQb0obW7Sxh4eyvcDMy36m8LT1sCtJTbt11mcn5BHqDc+19mCFwL
X6YMzGdhJglujBz1ODMyoPxBVbs77xYixzDFJwCVaeIo+j21EiWUK0S42UfbTXAAt8Vv99CiH2GD
s13ZqfwhIdJf5weao4oXYvsn0luo3zuPHjfvINgc5O6i5To+CLWIKCPd937jKadKQrTgqRBizY/P
6AvF90NL06M4dgGZs2J558E+FMTYnqYh//fQYc1KGRZnGKuI7f+XwACKRdzoZR3Ib8+TiIPvDENx
aaUOXLEzpFdVcVE/YJtPG10PjJHsS6Sj6usQIcisVrhfJ00FfUaQZs4EYt5mvDclm8Hi+YlCrY1L
qTQ6aV3q9mlL0w2cs4RV1FPzccS4E1tiFgKelFEQin3I9mUwIVYWK3aMUweJiwZbnhT+N2yKHpQK
BAt4UQiZ7z1WlaPfk6poq5MKh8FSlvpH78/u0DYUC9w9lGqt7vIeAsebOnfQnOIpoEXAMlKmlzim
8v+bXBocuaMX5XYp/YetXCUlF4FKE7/EAQ7iK90G2dxFe0xoPbUrL3ctDW/pu2Bb9QxWLsAQlWGZ
880PocHNhF5yMZvhKQnfIvZFxLenLTCcdnXXNz4HWjxLaeb+PURwMmmG4rT5A1baICzItKJy6evz
dbwhWqeF2WkXPA8RcRa7hMA+SDf2u4q+/1nufcsR9k0yfAlKHWn7a0NFFBIQm8QcZNdvy59iSdfF
xPgbS0zBTEhVPDmfszJATioJtsOilfHjwd7fSQsmW9wHdCx+UvO9E/VLQX/brueImKVS5+nlfOXC
NDYKCSzxqpHjlBGsp1Cfk0tuGo5QnvLe+/RRvAkPD8giIhHo3epS8szrgL66j28wSXz93pa6+w65
oiJgWzmp+5WiJUEa1j1agfWZfUbr65nAr9lPEtzE/aGnZxoxMCQ0rD/ZwUIjJkEqRdvmbsGvBbnZ
X5LKXWCsiKY2Tc2P/sGfN85FGcGruyGYrXZfscGkxaha60y4GIJi8uoCoiF5fc+X7jv4oPNxr395
/cKslH90VIHt7969FKetCu5FwNtRQEI7tAuxGd7JaFTYfM/s7doOyWZ2rJNbdRFLHWrxgFkimtbh
3bSrv3XOSNXoPgIze8HO7HIancIOK14VEsgA4WUnPoIqsNKZdOoVtk7fpamAZB2VwGq6GLY6yO7P
UgeJRRdKpB8bkuGiTi6w4JNC06076a4G1MuqOs5ohLQJtz0XqkbTCo/NO+QNnyv0aHghgTshmg30
uIcyZA1MThCb3hJtdb6++nZNtOA99ec85sGxE8Lh4AbNGzOEMtNMGlHa2sJ4VZL3MnvO7ElQqa+5
V4uv/w3B53S4nH7Ay2NM0vF1kDXe3B/v+FUkx5ixrMk6i8HiVGnGtk0Co6Smzbr09B4Ek9Vp7N0u
M+/m8s+ufM4CGAUxL9xYcW7iX+1L7PMFu9kEC64eltQA7/I3JoZ7JyrDJba+ZrqoBXrf0BWT1Y7N
sh2ORTmlMVZou7RMXiV+DvsuuPg3NKqQ4+MJGcBhcnD7H/259scvt8jLtHLdRgE+EPSuXMobb7pk
uJGHv4PBbz2+NFN3MBl4lB5nDOWLn5mqyugBwoe4JfezbBzNsRGeTetjx0bIGZ1lb4rZvGVj0V6N
wmDSHTG8ZM0y23gYchQ4lwLmHsmRtB0bwXJPWdt17/GjjoGOF/YWvL2ULAHI1Oeqg3yQd9rU0mhP
9iGTt5JazeuTcWucaL6bPOTMv/OXfUACF8kYglh7TDhMFZNihuy4dmW1dkYb3x6FCmfKVsSSf2R/
SMVvRrBLyxfU6NvWjAbq9MYh5htmEdvAE1oW1VjkQR3WF4R0AuWZk7wosiBpGi6zjiq0D+Ecy8E/
nnVIjv/dVFXPIrwIXpVU8fjdLjrNeU1YGpnDb/j4PIg5xothWyf9V2HpkLXDUHoOk7cQkxF/cQe5
uAdJ4FBr6doGQnb6hTqtjYrVN4aUEUWtmnHoVYWXz2QtOpJO3P65H3OchvnN2xy/x3VqQZ5Su6PK
tefQLMmZkg932m/ZDIZOCxnTm2lG1jSAHcOSIoewUIjugl3AvTLgNXD0+yqU3vydPWd05MvMYwe+
8a1db6rW23x2XL/jUDHnE0iuh6pPv6n2oXUkuRCjYHjMMMgSSlShBZ/4pPbGNZL1SznvURQE/30b
nBWmogqB/UJ4gxc4StFyCfv8wsQC79cCKXSdt4W9mVTdpa6yqI9jRvBcwR6Q+8Ccq7WQ00Hg0+SS
YIvql5ijpZF6zzTuVBKCvapvz2NhOnPQueWRgezlq9Yc4y4L98b8F4YkNy2CPvHUTcuIiufe3e7E
U+vZT61wun7hcYe8OvpaJDChxMpGI0NZl0joQiH1tZIp5kjNXIQdHf8j54zIH4SnzUKTcxAI5kW5
PdmtpDkxkGJVziwL/PUkm4ce+GwPaQbCm8p3ELdDylqWIhl3NY92RgpUB9esC3kHbvcCmcUpxjpr
/GTVhBaPpQw8Dy+ylUIM3IaU6LR8Ut1XcEXF5T9JOe79r1IhedQpq2aLr/nzX8jLoJRq3KmwRSHY
V9/pKMumg5fQeqoJDT0HOudReDdmA1ymwWDhHcvfiJFb9HJJ4JEpUS+tXI/NsRLe6c7mjfUn1LZe
oliGsJMbrFnHBbkAI9YnWzBe539TxUsqvqVVil6ccGPXSLp5M+Mb0rknJ6xfN9cexa40iEw1zFI6
XCPt5ew8vTF7tX5uSq5ZPG9gi+2x6SsY7RR8fpIWn4/JIc5LLDlo+NeUDR8bfL+Xhllb9l6weP9W
tfBZUy/lASyHy+NxKWdvL4nVKJRt/rAh43Z0VvdpBADXRuZeRkjAcslByDbyOixkrLoFcq4tGL/D
7m5u278T7X1HvjigwAEA+sjgGT7vEbBeeZzZaf+YAoN+hmgEak3vkImbebFlMmR43J2uvztDAq1i
M3BS3ZVd3+8E6G+5ZeGpfKiMEAEVq13l98I7niLPDao4tejhAkKxeViojybONvQwlnYJJ1HZFZJk
l1CYgQddx47umflLQfkOwRp7AmIo4L75DGvkZadnHzLPvEha7xbHdkVIZhZOeC96BJ2UJczehoTP
zFg7GNrJGXJ4R6O6QwNsyzjQuRgBswHAv7jX9HwIklbfPMBBq76D9kt3QF2Zj6KI399UkWzdYM/2
CqGLq9UDTV8TFHeD8IjwD3a1VqYg61J3w1zCTz8f5I5n6xl7IvBPFDk2hhOM7Rvuw/15/gNOwtKk
uRuGdvhKcLGUah9ihNz3xqhZRUv8Z9OmHXNWbksxbTY7VyQczSTq7v49pHFyijC94Kv7QnviUZEL
aeudhnlALpGvZkcs+qWPRT9IP5gU0NZUKUZFejQrhfo3J6+38gKQnCp4adpShuGcLdsZ9OVjwYBb
Mn11njP1vJatWpopgCIa2pKakde/maHfLO9+38QiCqZrDg2fty6QOxct1zXk8gFdJTCW2rerqh73
JY7F+YleB1vj3MX8B2HaBNBQPgdRs2hwlP6QRSmbQihNw55Etm47fq9I72H4o3LnIab2e7w3hG8n
UyVEKN7qXMCVSPOijhxnnz5JVmTI56I1aFcQbgd+ouuw8wtgWv3GtuFgpK/SPKfjFh+4q05UOcfT
Tl/66d2q8ZDdXLybeeulOUV1ikHzVp9Jx2aPQs9ru6HQZ9uxlcY8aCDEsgrwfoHAr+y6Z10miOVX
x/ewaG5kjEv07Cl5crwSBNXnfZl9HTa03jRVu4EI9pkBo2KxNdcBdkcL2KoKmpYpnoXXPGRdi0eZ
vshozgU56wtX9FhbzMp0JWeRH3wCPh/FyZAKUKzW2IrWdhgPtkWSmdoqyTPweR1fbYIBZ3no/UpO
OVzSyswCjyGmOGKuKmF1DYPeYp2TCw2wrmtsfiGQvYLOjWC391T/X83ldWt692EMbVltnUi5qbMN
VU94j49zO+xN+gGBl0m8mjhdKzrRyVj+kexNqwSG72UQY5aN6Uzt+oEjN5y8IBAR4dB+R/kpXz0Q
ag5fi00zTDqL21hM9b7eG+RLe2buFRUJj35WgU45mbuAwgF/IhEGCFpeEBvLq1xnwU9x+LLXvZVY
O+9IIZA1j4oqe5TiUPu4pyVhlN2XTAfCbYd/O9tlOMQxfJtmL8hTy5CwS4w6/gRLYo93jXDwcx7O
Y950ty3jn7StI+8FhXUf9D7AaaUig9fwXzLWeiPtQXE046bK8Sx3zrI/ItX/p1UgiHP5dyR0Q4pC
aABNgnIg9hOiQ15srQy6aVQJoPFUdsgWzbTTxCUZlwSo1XT2fyAOzxcsChamMH+pAR/5QvTMmNQQ
FaaWgNMsI/fWP9tPwjQU5CsjHXY9LgU2PD+BD/ZFzq0WwMBFfLPw3Ewk8qiZjG//Exg5C2u30D1k
ffc/QR0mXvCyHL1XZ0vNv3wVaOrnHQIyVuvv3LIVxI4DbvSb2xbRWbEDFzngqfVox7Ysjf6Lvblh
AAK9s4m+s3c5UO+AXpvYJQQRq/U/6t+tl1RYFzpjgMcIqYUZJkKeL7ir0Sv46SH1Ubqopwsla2jW
UkuQ4o18nn2G1o75dvdygUDI5Bc3QXhiuWxYVHZ5cqC2AGvjz3wfsNRPEazhybs7oNOd5y+y5HIc
R2KaO19jqbu3HUu9TFOzHpmv5dU+bYhgUWWzUkhdkZbaS2jYDLqmqBylhzlgeL3nqKV1JQv6eXFq
jj9zqmpT9gN/0JdwzOfRlmaBbk2xJpdIYpa+NH60VwZix8/3LDJVgwVXIi1+AKlY/KQd3vp9ZIaN
PmswvB1aC6PxKFgmnBENUP6TnwYBkoxJfWFeNc+3KSTZJ0tk92FwS9X8FttDHtKaGARDt+ww+Hb+
WpSvTpEoc5pb+ltKFK38Qg9Y2lLx1FVUbixVEprxvapxmf4Brqk4a1FRvNF7bGjryFzw3PRI7Ffn
xiETUCnV2lbDXM4mp9qJHxCO0eH4jSSf3Hdz5rtKir9qXwAnG0XtWIIxGSt3exRc3lKpYToi0Pe3
WsKwP4UDt2NztV+OMaY7er8ik8Ey9C8eGAQMTJLuvFdGu7KxJ3dCaDXJuu5hM3J82OnPPiY6JVC9
Zub/k1lc299ibIACtH5+RnYZ7GYokwcuPvXXoZ3M8RagrTOlyTLnn9oLIrdFgNXhxv9rolocBILH
bQzCDzr8RIEas4RNRC0K5HKTpHmmm8SJ2LALK0Lu/qm53O0/rjArPtcYs/KiuhntcEScBjl/SA9C
pPgclgrMxcOLu0QCGGX0isqmkQPkbYevhdUr5FPG56fV4vt96lmARwTRWt0dumEM1aqsg2mGsV27
znCD5thps3k/d3isVqQZGPdUEl/x8vA4BNvy7DC6fZounAppulX7cbzjnfWxOZBa2TBiuv8y4G3t
LsELcjSSDMYf/vS3GoNqVi3wBLUyoqA7X3vq8UZzyfU/6cPfj85Gs+d3QVKFost0Vfn3An80de/q
zUhW7buU+P8OCBw+eoWXBGUAz7dpVvHbUFa2HVkXwkvK4J4JDYFfKBq2VNi83JYFZGTGo+WmMIbm
G1BCRhrYv+8jK6rE8mgP9L3SLyQviExjdAcirRd2HuYj+yu1Up60IJG9ER0x840dFHe5eP2ctHQS
IIcNhts0w1UpQ9qbOqckBoTkPSpZciBqWvZGVzSZCOKTDFjJ8z3kMB3Amz2R/HZcEBuLEPI+qe3m
GDYik3xd9JD82LwhE1UBc1EtpiPawXykmmj+j+dVk918vQjuVHDKdFooBNZXgTOg8/JgkRZTS6gA
9SNVp1GdvbabF/Gu5XJp/0tDGyY3KdiwRufAsbADATCkLH7rFTjPs7wcyfpz19RlVxHOX8lxh2z6
N4/bWxCvkkdMvehYoV0DGlhK1cuvirTef4V5nMTta0JWwbmYIi6glngiNvR4jkD4i3Ix9/sP28xo
+xZeAELRg2Ty4UdH8CO9r0VMOHBoPFtqClatVceNTgmZKQ9KTAZ0R+Fu+00bEGleEsnEksBr8icl
UHet5Q63A9l9egWLQTMAsoAH6hoFTvMnNzl69LwWp/uyaDBPzHPyl3Vjq8lxLTZhFa0l+pKOiIAv
ZvHha5/hkD6VddEf6UPU97shbt8T1cP/Ss/THjwnQ7Crq+SNBWQCKn1xPNXmdPOYCW3juy2XB0SO
4erTS8mt22bcuY0vPJ1e7P+YbyHM9OrUnan1pkPOEzBl/aj2N51IMwIA1aFPDoR7v2osPZvdxTIF
gibHUGnE2uQ6u+Rz9yY8KqXys8jDjq+XpDY7AHTd5071l8xd3HP050zC+2RYX8IbWMAajN7V9ClM
lmDMEqKvG/x5YWKssQAtXS1eBw8FVb5TAo6u3B5ANREA56Ao+Bg9wyBxenT7d+kMrbrRMs8VL1GW
/CtYxm3Zeo72Q+mh9UgYasbS3R5BCT+U5GXQA1/08Ty8fAiO0eOnKBZFjBnx7e1iLRFah6wXCKY9
SuP064W5m7sw73UrLxDSw+Xcg/5hz59w0oBSNsJpM8JZTWGe8R+VAkX1QpAORHC7DuAh0XKsre27
Xq5WLxcSJsjnDclZk+usBBSrU7pz+dP8Dvaq8l44IEmzy/50aTrf6Vm0QI+L7AdCdX+EYWtOFHEJ
vph5Rl9sGa1zeITYDBcMTT80adtBBhhPAlxacmtXEFL972BXec6VSqciEFGvH02/skOqK36wpAq4
FmLTROtBWj/r8SuxVakfzYtny29xlaQ6hoTOZikVfNY5L0N5ZC8v9dG/5mZMY13XJtRZuxqF2umh
RMrMGphycf0YzmmkW2E0ZZPic0t0cSnL3e63537ZYJVGTtFuYlIQg5EVS6hFrwKVqtN6KJSlcldQ
ueawD048fJ3PtPHsrHce4Uys/b8NgbGcFlQw0ahsExWiREGI09Wp9w+u1Alyjw8Fb1wIZVurPsmJ
HwTUN5VsFnUemOhfTd6RBDnXH6Q5RvWadXs50TMFnMMPz41gUhq2VVjDB2IDKMoHOeTQfww4sTkn
/6aSroLptnRlpPqM6onEAtcWTnddy9tRpxaI+4W4gN4C4bSY4zZxKiF64wiGSOszpmGa5JDGyhGO
VeWUxwFM9K6wbRGx4ZL9fLEf5WFa2HhHQwWoVuYvZRFmvADgulBonDVMYNSj9H01S0lQvkmtJzss
eUudVCnNF/wFOyIxHU/nsfaDlQllXd0AZnV45YGnCn8b94C3eFJOmbCKKxBCAPuZuldTBBkUkSWo
9P/6fsDRHoVWpiD523A0v0r5oT8rL7uGV5z5xZ/zsoVCHkkLwPkBkbMd8DTBt2E86sh6sNXnlho4
nmePEX1phOlztL53yEicSA/uzPd3QX97WWbQZz3F3zoTTObUBSR1Gc8hqQ9BTLUeCza8flXZ8eg1
dBWomSYnt41IUR9tDyiDPZim41mjmk/y79CbYiGlVhu0/ke+Z9AvnwYtnDwBreMMFAF9YcqKKL1O
S/uSw1zUM49gpEN0e5nw7DSw1WuTXfYoGRtOTlOdVhm3nUmeoDFUSTkIDU52ySZh/VpFVgAENc+m
Qa6jgvrPh1uVATGAoAO9vsnnUcnEHWwN3NjWrtQXvA6tRcheniMoCfoAdJfMqH3vxC2bvPhFVAdI
7TaQGO3Mz913RgMpQJxVlB0Hu2sVdx8WgwXe2/Jlegi1cX89UOHczq/5afyHnNFE/2vEe3hGDCBV
4FwKrKmdmbhRrWUfzmlw3slSoEWIB5GFx2BuulfP62DJJnugDDYDw9DPFht+C3WOLSSGhkfvh9AZ
BL+dERDUV9bT3yUIOVw5zoUmB4zXrZ8pg76LTrRGrw8+5+peT0TEQWexXXj0gVZ/Iw+InsW3HBdj
ng+ADVl/feoIMryuyMHdtBuNQrlKDsEpqxlY9MkvpfOSL02ppJQ4VZRPigtT/Msruu1kDC/dadCH
xJpJb1oSD1WLTCtKa6zHxNnzB8WtyvTLEGxsw2IkKBeFLzkTsyqQi+UasHgsvFj6LRf3QvqLJSN8
4DIGThk+H8SHtWhedSy8lmVBpIIDQViKgMePSCLNT602OeM5rY3J2l5rbQxgt2M0ihOFSDP34oWi
UdiSdjrctQLG3wIIMY3B0jNNosq44/PCOXZlJirEqh5hOlrpkv5MDxb9+Qmcxl7ZW41rprY9crYb
3FbSkEwYtVpWNGL5BEySQpapEeBeHYJ7cL0DWpo9hfDkwBdmIRJnF5HY5IQT64vjo60+kQCpIcom
pgOYT9CfARzxUPgMulOjP189bJjzsXPaPVqNupb8tGo6GyH7Li6PcseqWXo52m/AZ2WG/s4mxfev
mHTLi/Qsy6ZP37w50jp0fU0hnpyIFptvfLCqvefqdM5BmuiQnj+fvE2N0O/9fhXJw6Q3AEJ+uPSX
kkAZeLyMV0VrH0EQGNNFE53Kp2OfBqon4jpVqmO4hpyi9XAg5fUtT9YJ4eKLYv8NrXDN3oAYa9sJ
nhAnOByABh2akIefieS4EY5YfaUjbNtvytZiInSZgtkAq8I9ip3Hi+sGU2Aasr81j0jEvJTmYMV8
Jh38urOK9nrlLEMPZsyxJm8ThjM8/3Mc5rhAQnV8wvyiQS6CSUy3roVvBN4vCJ4RNIkuUPnc8W49
7CiAKAvTRwgqw0H8gxt/XiDDbGhy2sPS1X1M6gd3uHKdtrdH1e/qgj5HRE/iHZj0DWFUD2N1lGJG
pb8QLzjq9xBRoiEkwLy/x6kdRkH+++GS2CXitIWllkxEKFMr9lApVx4ng48IBPrtSfN4FSJoGI1P
ROhV5OxU4ZMfsQGjMbAxLBJlXK5+wnGeyjVzrHjO8+QBQ0NriToKD2XQurOBEVQQdxtzmwAG5aqA
+FNxyUaDgJHEtO8QsJbUwl2WX0gQvxAhmP8WHdqjsTEBDhZUbevHwd85OcHWjI7b/y4XWQx8R6WP
dYAX4ygJM+PSc8zslwwK9LEDySxxeUpf47vjFohZ4huLTJOSHQwCIqwDlGqY2ncDD+Lwa2R2j1o7
F0gMBvWfWXNwhF/C5uob4yo/kXJ4SP7LcXyknu27KCr/nDdANCgcqRzQRyyP2y2OBKLKTgR8MZvc
57yFwBIGsJEmR2DycpS854BUIZ4mZEFVE/dIB3uGa06E2ECGoPVL7Sj27i/ZdszLvtZzzRk3qjfi
WsBPcohdTC9hTBB8LD9kP+4TE5ZwvzEqAHyyb0jUNroTebCUwJ0Xx9MzRwauMfdyP3bQoSiIZJ4a
C4OE3tpIvP654/7QWTCiY0UMk8QBnMp+lHYPb4RZ22yjX5l0pa0sVLIq47ODBcJJG4tH/DK+f+um
hpP9wyZlpyRmkTJglXWpy+dc5WIGX0CQ6GlJuiXYBgO+D8TvSR7VfAGc0L5uHA2YNMuktMesSXzJ
NIvo09zBxcwDARwidPw1LDogHFXl813j60znd4SWKuRNcUHDiYz8xXU6qFW7s3p2S2P+J7guelRL
tPNxvtyyrCPCHjbHPQjKZF7V7RfgDf77B71PGbnKBcoGAwtUHn1BGF6RFjkmgUafhltgiY0jx/0U
N+CjRZt71QmWsTVsIjvqCRidmQFAqI2433kSOPWyxhn52XmfckmDfM0kkt4bpJVZhkyPYCKPWLtp
bhQ23NVUkFrcvDJAH105yz1FOGtgVH62DyoecKBNAkOsg3I6UWn01dnnBB9U3PltmE9+oaabCyA+
Hww3ddp8embU7bS1cHpmjzdNV+djPQHmO5pm5mI6uoFG4THGpohbbnatdMIph2DUQBQyU34L13Mr
ueMzik70G6pRxcqmABtrVkjzYLEj59PffEaPi2nKPHLB2ehmJ86SFhZ5jiEd7Qx55NIH2QC1MuDv
CBaGAPkDYVmAcLe7jKL8Ai2hTgcfjzILaDA2zCM4es0jGONmtPHATSu/VxXU/+IDMUqdKjVLL+00
0xalpZLwLpjxMZAoNs/OdjwO/+U2Uc0xtcsYj2M2lM/AHd5Fk4T4YDpQxUEnsbWLYOgol2pKkWTO
Bho2A+zTc86MX+SgUweFEDjikQVxJ2D4HAuQkkbhFQXcV434XxWOoOUIHzjkAZDjTwB5ONdOHQ83
H40dTAgHyyC3g2vEwfJtCWXCFNJlT3Hq1KOTeebjQDghZTZn9g49Z9Ge7aE2Bz9eHyG/m5acd7KP
hFM+KrWDzdbfi/JpEkL2ZDbPaQE93Ygmz8toIUJ+3z2Sb3xVEDhWUmJy1jz9DJl1raD9uLCu9Lqj
UR+hQDCJ7JNYWvHdD/FYbyTOmEy/M0ONKz5xAj86A7UVwY3avOwbT3OOemXxSpLdLTpcjzDoqisw
4jsN6hhEL5H4Zzw7IirKvW7L8fN20qCdaydpnBBSCdYefYwEgU15TW0NX/1swsG4+tnD2VDl9jm4
8HQfB5bed1r1Oyz2X9G14jmE4yybeWHaOqdRkTsxexYQMmoylh0Q36cu4MUksVTwTIIaQqFu5hZv
ck1pDjvLcdhut/MYNYDf4YoE+AWFUAgMaaFvTIbAGbKyrziLvWhzYqjpOlBNasxLAwT4SmwzsdaC
HLzIb8vtE3JWo2Zk+w09loHRwP3ZOU7cjEg+HnMrry3EbhEAfdNNPfQj77G3yP73yCwUNO7/CuNs
cVQGO41CHR8FwtNboxqDf8Tx1sNizak39gZIHtL45YADYat1EUPkBa5xqSmhNYaNbKVVRv+RgDze
txT4mQUfMMQ86SikTOShuZbSf/Ou4+x/PvUWbvWnqkLGQSGdpCSlxSD3K7yKuKK0mIHg1xnEdKhs
y0vVVFHhQzjCJPe1KnQs+INVXn2BqrcVt4CLpZMv2ZpMJhs9t/zJNqtCnbjLHBhb9V8oQI5t1dcz
5rlF4mSttbd1hl3OS6+C35RsZ6Bg6rvzoqhr7AOizyZQbDorEzFfjaD8U3RyAao7FRtXGihEZHz9
CKDNfx0mmQqgpktwbfHe9+wZT8HKB+MdlOCi1c/isFRuRr1PsbvWotJK8PFMnV8H8TI/GjGwu79w
y3Iu6QD1YsQLO5HimhjuHmwAEeNUpKUKFkOydE+2zAdjZszIoIRg2zM1DNUW9AbEwSGcUEPSSTks
pjkh6zHgbKl1PjiVcs+IQ2ABqYmgvHegZTJvTt5WGkk98B9sAoXaPeJ7AuvVqHFrtMPy5FP4ld0k
zMM51tMyR7V/UB2JGvch+q98YJGZ3iGvgbLV7L1tBgEv4R/NiEYgvjqh8NbDPoR+tuHmyJ9StPw+
GohOUakU7hDnAuKOQ4CBaIqzT1+xZwnjL0aGoWO/TQJBsIODgbbBmmLVEMGXkR8DEgxCF4kx4ulW
LWTmFe2XjSSJAzy8lBV53tvYfGZsSfIeA+OvqsdtGxKCOC7AOio/qgr6aSCdmV0m9ue/YwDXK3/v
fLdJZyd6mZFiwi7WTYjEShb5HxuU6BHU/F+8jvmQSin5FWd8XJkgftX5T+SzmZP84dkkArWRPsSn
mQ71XWGavr+yOQFPszuUoqIpVL+hrDnTpf1dkVoxalcH4D8YtJYoW8n2qgIg/2CyTpZ6VE3uDu9N
3ULzoh+IML92yaN7E29OFaZPYs4+RXkvc+WIRR/OvTfZT7Y0f1bprLBFeU3P96wudbuz4QvARVOY
7tDPU2z8JxbZoA7INnTIxwlNtyKe8SdDa+/C5kiRUwlgfG+Q/EZKek+LgB6HoLYP49g6Lnzde3Xq
AEHj7DijsL+FBlt3sgsvWe4j1/ZNq4eeK+aXlOS/PbIWcv2YGxRb4aRNS0IfhMtQLnnjY9P2Yt8Z
uQFJG5hhNqBjwYh3rDlfIn2MdpPJ7nYx+agA9UdN6hU2SVODfZQqLdTIkEg+iBdyP/iU+p4EQsh0
ZIGjujFiNxKpJBhyatll4mJPXCRG9IErKQS5YzxEo09VHIr+s2tCylGEDRi3nSsrDe6azOD8pjQe
wSPTPGl1rRtrC/AUTBIsCkDLsMpAM0kyOsspBDxK4xAF0Or9LkT8S3Z00EYdSq6RaLsM/5msz94b
kQnCas/FN1zTXM0ozSeBUZyc448NV9fvrbinbUWlUey/MGIoe+yOA2VpaLw4tGWBFxNKUQ7WHs2n
Ctt1mJ4KyJt88INGFK2kdZUVh99PAC5IxoJa1GmOcHmqzreQvRSt7dGo0deNmbjpHDmCUwheHIHx
sgSAXxmSe022wJAu4dD7u9YrGQt3Qpy5vDVRrcT7A6goCvBpCHsCqT5FD5AJSiBhRoyrGbWzU8fP
FSKAxpaxAEWBoyWGljlSMfWwvJlDKm7AKFwrslGSN1z0bwe5Y8eHIhA20HRwABMFUkN90rNQRQNr
0r5jx3I7dnCIMAm5sA9DNrOtMf0f03+zBP5Rnr3gTUsuA4vj1cJv7o52FnqgchtgnUeuxFRB5iNA
cN5egP/iS9PshlpMRB/W9gwtKAGLkcPHmhLBk5nw4BjmHdbFy/7/U+80E8tRIsJ1aTLwQdpHuHJC
3e28HyxVsiVOHN4ThiU9QF//5I9uHZrVgPeqOSk8xdpJugqXWfR1zg7RkCz8b7n209K68+0Abemr
igAj9156gd3GXYpofm8fo4BUcw9xHQTZ2Qk0lzMj2bpfcN3TZQjT11b/KXWMOVtpAr+43KG1uhRg
gD/ZVWqqRV28X3oG4ufSH+6sRe3ji2j6WK5jO1YCk76zpzfFGZvIePo/Ib7fjtvnhoilbU8dvyXw
CNTl166yCGRkFad9bXIgEQmKuqgEs3SFc7gIjNK86KEaVdyTobPGl1rj8pHLClrpGFq0Fhkq6Gx4
7XA36DQBtHiHTF+Vx9zPbVd8SxMapIxIFhoP6wLe/WK0/Zmrhc7bZjuUDNP9M4+F8l4/g3RuXEvH
NNkFiDiTI8Rdz79Iy06Xw6fmnE8X3oYSqSty7vUeD3kgslgmQV76vjTegk/77lf6HiQ9lxjnIQvQ
MBsjN9PvIKXNSuBpoTEkaT92/PxjDxFU6Gtihw8+WMhYbCh4qIFxABeiD8YSV2hLlm78M1ZrPPFu
s9hz3PJVODDq4u/IdpTve9vhzKtLsZjnioow6ZL8sS6AKH6Nqo+QKHIeWVVhYUQ+FLxLoRMGyG6c
L0kFF2PYzvOHfxXYh9QY6K/452AQpxgoXLTOvLjvVyh+etzKS6Bl3BanC3cXMPX/UDZHLAFZDyOc
qkPQTp+kdUejqwoGtbqxCO4PiaOtHXnRYGPkDnwuV4orAxbbqFv85M2FMm5wB8g9BjmDAdJrh93W
MMLtb33O8ZsZfx5wQODhHcuncgAPkjxmAvUpz8m2evAa/7xqWPtXxTz3KCXoylYyZkH95GjvOAdH
9u7oOUYBpPWC84FxJlpB3i4KRGJ0Rsk5zQD5/tSPbEVlboGju9sDo5nncPC4/ItgeVhi/xzh7rlR
qa3AyNybpsL5KTYqQmw85RbvLdydjDl/QbIdIJkVSi3lf4BtFWbHHfjSCRIhGR8XQwPIDZ+ovvfn
ey7FErpGoim1HeX5VpJ8lgW+8I6hQCwEHV2/65u43htOmFXbLcizx5MUZVeR6kkkft4mff4mMMPv
QmrFJA+ibweSI1+/ec3iSIHd/EtseSJQyoaYwLthNzVkjzlOz1gwphMXoQEO8V+0xh+ZwKdhsitk
5GMwTsESfocaCG6lb/RVL6/7CaaxdGMIAPxfn09IUn8h6g2M80Lrv+RsUXcWhp+5GoyQa+9bAuee
OkNVG2BnwE9V3cscbZy3CpIaECV+PpMPEck8mqUYQKtObtKUQwm6iJV/msEMBi2hxVmt54nGcyNY
56njZ/JloCHpSpMzP5GOPa3wzU8gbwdIWbw26WuCkZ51gdbZve/flFjytUt26kKHG2gDqD3/Qodq
oSQf2FEWcp0uZd17MI3dxDT8X0v0pswjNslr9LZ9O0MoOgp6VSMtG+ke84qcFf6tVy4OgYPa81lF
O8jTwwPtJfPJzRT/jJ+1cvNz55t1/akM6Xn60aZk7U4hOXH7VfSEUuECFJLIOmaHywUzTpOn21Pl
iE8LuLzrimBmZ/w9PAw48UIe6vLFEU+js6G7snZiBtfzICxoPaeGgypIMpqBiBRN23vPrdh1JIb7
FHUVvixHSfen2wT8xCb09a3sXU1Dpisyj+Q+m1CPKQ6NyNOPluhhWNzbF1Psfhi4Uym0eMYMwRqH
/iizIqF7nsxrIMnE1/ja6aqDzKeCU/gaNbvTLUyiHG0PX0bflNDCwgcFnbhJdp3Cfr8BK8Jx+F+q
8Z75h75cG4qFd0GrNO3w9/xzqRB5W0/lNy97cHW4V//V3vk0o8H0Pv6KBkL942QaCk2NbmdyRReO
RSAXHuHh/LoY6166a42nkau7ecy++XLAMqJvhjBUA8Ebv9xcZwzYIRuMvcvbMGGQYHiW2/iIkEBA
UKkYWlyeN8tMku9MFKrpR2yPlLArM3b+i2qTBYCzWE7CGrQ7jQscLQuzYoe2lODPCsZYEnh9fr7J
yEJ8+ELTpraB0RwV80XzhFHIedcdFtFsbrXSK3hZh6yCVW/HV4NWpoEaDEizFdd6mGcv1x/5B0rw
TuCKSiwbDfPyxaamjVGhqLdAdPDNU26CQnC19Y0PsRmL/ZmzUfWrY5hmU9vPBUnnRWTTkYlgFYv3
7Y3EPCliy3F2d4UdNLPQs7L5A56HNgMvnVEUR4ogiczpnFywPqbK/LV9+cVwQQE0nN+AVU7umcQH
e6SoixO9pM5mjARzWVcfjW6Y5arcBewS7symbNYWouG0Nc0Co9qUoPmcqNhxqg3vpMWVsEeAVEXb
LiMcgtG3/JjyNglh18Bl7tyh6ZjpL9epMzuxS/nv7PjLfvc8GnNG6kRDcZ4rvNG7M+jYLaV1sOEr
XBiy4lq1nqlM9LUmKIcmDlk/TLKdYlop0D27q2GD8sh0KVGbvgGai0x8dv2w3icUquUVizQHFaAJ
W/M0rhyHX63GYosoUfyP8MndU3K/AedgvBn/DhOOoH4exhsE7Vksgo4XM06KQz/LuuywHgtCrcIN
yg5OP7RHxDBa7Z68qcYWxNG4z+53RxqenaK+y8+zCDdL7JKPtSXLT3/Fy2gxY4vbTZa2KQfqd09B
/QDX0xiC+5abt4PWj2fD15O17gac3eVlHo5JqW4UOkfkD30UoQ0gwVhEbP4JdPHqaysecs/zy/Wd
QLTvC7vY/d/LI3380IkoINFK+oKFWzzAcRvD7aom2tvNjMf2enjFoVo58d/UZR8dJ08YvkuzHjyT
uHyzj/N0fWOKRHymUC8B67S78IwoaC2I7d7IFvBGSWpkjznJTV+z0Iyha3uGwVk3+eQamjWFzgUl
Guay1RcTVu1MgGtQqehG8pe4Gneew5WApm5FExMHZmDFb0Rjxm/DzpF8XY7hXMF3XBw6TL75zepo
iKyRwGjHjc96o5QzKcsiFO34KdtJiWffjPDhjClhH92LJW5+20gCURSYXD230lJmsw5vxHa5BFWZ
poqYFFmksc46gzDrFZ6hYKWIFyIwzxHfEnUfBAJBzh3mHTcl8GfabgSAi1guM4T9Oj4xKcWKkVz5
PWaDsejHevvi/VbsL45LnRWiro5I0E7ItadTT0qD8pBNLpXhp+Qos++SvSJBt1k5ZsPNwvh9E1J9
w5YSdXzG3VAI7/bDv3oGUEMqkFby2ajsLEko/qPLp/gl/12HV/UYKpCYgIbrf+PedRryPD7jicZu
88MKvHd78mxQm2aK08LOJ1Yzp+j/2fgJUXO8LBKprQo7apKmkArYd900n4Lu59n9K2QFUaIIXc+6
ZF9L5IsmHTO5JZHX19FXKDfmfvFaCCyhmBxlTF5urgLk73rh1TtuITTRvyYQgDj2kpWeM0wumPKy
IKXrVIJwPIGPVO+i55NKklK7TIqn8Uiz1Hb4sNuf+eVazAMtVoM9lvII2EGakRQK77RcluVSXM8p
IS7PKu7gZ7r4jKM4sy0i0Xa8csMYQynMMOgskioLN+c0ZTz817Z5tap/RFw2VK+vaU6dSeK35LzU
ozXE8P2NItlu5D3Nl3fnjef3pG7dHA9tpIoG9DLNulcRJAocnj82XWUeIzFbOTmBWAf/wKcdV4sv
TwDUlEC3I62UNRApRb9QptRnzAyWhXSbizWWhIvEHpTuoO3VnNoJH/EBitvV9QYPovrepLhC9Xyi
suYXoipnb7EtPhloSUWTHnWGmkmhk5dajmFc27D8o+o/XVIVTMLF8aqIRH9qKG1gBzabYXCTupyt
j4NW3w1fv5rljPaT8I8+sYuKtP+HdwRPD3jwH0ERsWWyRTuzKDWCRpE2plIRT/EiiDrDEGr0K5Y9
L+UK/153FCxnCHmRV9Z+VHWPArO4Duhkt3iXWm7Zk+tU7bT9edQd9Ww6RLl8O1XbYpBePOmSrlec
oh0bGw2YoAKBBexbkSSAANt8RVkQ3euZtbWzyOyEAUeSeKYawXC79BT1ZfzZkenMduohNi3nYFlB
GP8DygMAWA21v1CHlpiUgPrJ1BO7S8TGZZSSZDGvMkXfP7buyKovadjgmjmT32Vv0o3dZriH5zVP
QzThf33MjWR6ixBvJ3lfBPer0OBIDPuERradvkXR+t+h4WwE3cKZhNG7U562lRRYhHavjZOK5zNq
zE3kuqSwFyT1bVsRIwpazrfEUcq8XaCPY/cjhLByx4LXKrKR/5c++qC/tB3jgWGytI9zX5T3wKpd
0lHSlXPJ1wTq5hwnkOMXAJsM81lGbHJwqDk/o9m7Lrt5fON3iAcc/C7psp2jWkJSavnPZ3Us0V4/
OcfKt17svi1VkAikgeNC79luO6jp5bWU/36dP1pI3PU6K7hSVSO2i6BmHm2LQNdcAp/byybPvOal
1ofjRAoDR11KdeJlsxCZ+X0yeH+NrgXxCumR1U3K0RPRqb1jZVx1fMXAerMG+r8f3ayqtsp/zQrn
Ybx7FPk2oGv7fjnMmQnxIWvGiA+wHFyQy8CsPRvggxlj5kJ6D8O8dJW+tmmqpHcy/ETqgnDyfPhf
aEGuBFvOejsqKeIh5fmNueeocLiQdc3cNgo++4GtNuK0jHhQ7TsU4Rpr4SLPRcIispByqtxI4Dse
sODlqc0Q4FUHP4p6CgXC6jSiFjy6xVwjVGMu5XmXYIAftyaEiaN+nZ0fWKj58gOC7ERPAJHQs0NA
iIrL+PVT2MMjORVi+DY7KIHk1ua8nDImrvy6sWcU6wSg+zyMd8C0epIq0VWYDWBzmWRP0ApteGvQ
2+pgmPe6M0SDvr1tu2ZpsPyKliXdD3KQQNwcC4azII/o1bxhsSb+C8KK04fnr8wddR+gQYzuJ1kh
QJ1dllRspjicgZy3XC2lfzkPCH/2xd8EId9L+s0Z/8GeyLbtYd2XhPkj2TDqlTkEWZIXygOQJ1eS
4gc2+vURjzl4z1Lrl/Mmoe5jsalHxj+OJ6xbPMVG5JA1sg4M0EfkyB1qNmgGnaRQz8b3aohUCl/v
8qcWh4uFA4hd/gzgtII8j3NBVu3Zcgp3q7424eB2Q6daRXfocQI/DUm/7GjwiBUoZ7y4CqQ9ol/k
dVLoIJAqCJTZRZw6OUhhvgj2YI7RyFEXLJQHEhA0FxNfE0Fuix9BqMnlMDXZ0MDGgP24TbcieiQK
QN3QzJX9Il6c3YxF5yhZweqTZWWL8jW243Aff0/W9tn7U7BAIFSw9ZaV/VMR7H72+XhGYp+iVa3M
zHghxeSGFjTbGqd2PR+9KAHEbtQYFpPifAaJoQLtUhML5A2O++e0Ke1M1BOFAXPYEoj75Dzm6Cym
tWkavguCDACnD8avjTh0hFGI3Brcku2E3oO4mC5HW+gR4SMhm+i1XZQi5/T0t6fekKSmeNzZuxi8
CM9oc9wYgPgVxZDM1tBAYZ/KsJuz8vSlWW4B9SC782q1DlWRz/VFKVlUcALCWsPbL+G+tBoCfgew
sebIYXq6Q4Ncj7o8mYF9ETbCum+IGu4kZmoFQlN4ZvwlQIIsME7lF926/q4q45KxsIBWQA5lNl59
tcOifKW09eoDz0OfQ6UJX5VAN90P550OIq9wGUNAtm1FyRCaP7m+zTB5c7DtAwVDciXRKG+i5Q8W
d/qehk7yn23kXggvBCGZwc6Xkunc+Z9w5OsGZwSP+8jiu+/CV11Fdnps2eflldVdQeK9095aTuTW
sQfgq4xAdLOTsKnNtGTudxXyg5JERyNYdpe/nM9tefQOo94BE8Wn0uT7tkL9CJh9BLDGBzOapRc8
SOgZUcZyo+hqe4krLXZessw5xz8We5RsDWfb5rNTAp07zqtSNfPVeMQtQvWX6yqopyWE0NyAt8gn
A7s6P4huJECXmDn7DzTSKo3O90buurOYrY2bg51J1DaBtwxC77FSmBG7kJSZtF1oMdF9MRTevIrQ
G8hAvC3+WfMWi2C+/A5FSR7LuDQyrwDTfLOC7pUn9XlXxwdPd+tEP6tqYgDQ7DHvrPUgNqIkccWH
9rPW4qr7e8k72HJEo3dEYzjpNwmW2+hjOy1nsufjxkH/69wCuT3c2NnKI5So5xvepboHs/C22CzT
gpLkBe1lJfS2vGUMuRW3iofeHYyNVVm83Ecf2QFYQbbCxLZO+V4V3EItnQd1ELL1gP3q3mxCAqsm
LCmqJ/IpnojhkN4bjt2GpF3dyq9gv5GskSZIJtp+nVrLKsDjGfZCv6kRgOl9k9HBJ/2PHpR4JVmZ
E8omoAI6w04fGfG/aiUBrScM9eEqOX/6SZs54NeHZereQuOIVI7X9PE7/IuNIjP7y2ySnuDEb9U5
o+8TTzNvOzdUbiwVorc1GyoHT0qz27AbOwOJFZMfgK/EKoBQqHcPG00ZDpy7WaaVL4PrE9DFBIVL
L5CMNoAG/MhTPfyVuClqO8JC4cl01QSeZirPMoWmkG0Ac/IHGAbCmmX/5rL2reGjMuEmHoQbOMJf
FdBwZtnZdHIRVfL/bjV3JDl5fK/C7f6iaKwhdQRSqpspliZSLMt+knl8erTjsSjiHzOBlDcOcmWo
VS+VObPinf7e0E9+CQbI/iVTNvqrgpKuY+9yphEE92E8YyK9Vdygt0R64zfpyBBJQwHg/HgR1lVb
gA8b+FEupojUySE8++DZ3T064jOkCTlYxEkMjiyH3a7RCtxG7+xkT6SxgITrTBiOL2jMlmUa121e
2PJ26QJJaqAXJm5A2QyR1We6mVoipz7ET97rxOMY/M0MobdGpe550CyTJ1euaU2LwZfbbKQE72wS
OhqADaVsodCExdaioKbusKbpmjR86ZPRLfpS3/qfk2vaipmHHwi8sNHNgDJLwenH+OjIDVa6Tvld
h5igA/3lFKN2v2Dxe8Pn9RpcEZ5F09vbGLvUd0gHp7nUocK1uqtP3Tk0gQCJv877MAalbMmw6iKE
SAGMkt6C0kcxse1vN03yV0CdkrJ4mzJGPXE3NV5ZGUcM2rWVpEruN5Mvt6Bhk65v4l1ag00wCnLB
kQ+1ofJbiACV4DOAt1qvGuyjA8VEdNxbWJQ6ErXvqaNTAPLLwJBfEL99T7i8FHZ8GM6wa6pbYf8i
cAtmyN7J4SPsJyhMobkvFrYALy/iEcIGoZmjtHd+MYKTF0Kw10CGLhM/8HzgOTJeJqhiQMUzJdQG
XWJGLKqaQADJnSAnkBcTLvVFa6ou7si0hOWP51JnxZSUfkuM2YylvCDO9UhPzem+FLc4OfxKnMd1
YES+P3ocF7XNjZHv4OUjHp+zwUplQbKAo8Dcm4o8oh3v2xIMu6f36KmzkZ6PhVBtnXdayC3wNe9F
swDgHGchleuPEtBik9YD+HYm4iGVOaYYsMWU4Eigt/3ahpxdyNzrlZOTkqxFyIwp26vYlKQdXUv8
BtOfy3CezKfyXrDnLIDGmCDcZfYIEDAEC3ov4cKJYnTsXYL4m8lLlM5udPLpMGu5kraBJyEmfKM4
GYlOkwkYEH2YihCO
`protect end_protected
