

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m2u6houbd8w4XCxjJ7zyMdjRy/eKqe1WWlkQcAvTk+3gh6ALGcdZabPQ6z+0cNak68c7F93Hq0g9
c7cPsu2LGg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KuikBfmyhX0sWBVpqZE6TfpbCFdIEyJEtklBCeFBGGKD4buMZfD5oHElh9KvoFFVQRRn49X8p0R0
DtXowm1lzY+sS2gAHD2D6qV0gwFwt2GCgzRus/7q6jh+3kmhuSqaeKpJaq1dOCWpNXsFWSYAZsPN
Vj+PRlIXv9v2CiiO0uo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UlyjiIli3CpeY+RBfMdOTMCih1quPcfwYBLBz8d8sGlNOIVBh1S4IqA1uaf9lwS/h9sjnlT4GGfr
gwXBAanBplnhdvNyF7F97fZzdOVX4MmHjF8403wMjh8fkAdG2sQvVH0X1i7YlsmCbdOD6mpCxEbo
cyAUSl3EYb7Kx0pBENeeJHj0oV7YUnzxdVtqYxqs7xhyfmGSwrmrAc1Xrrm+oXCYw95RQZx29zAQ
zHT3iUVDHLItrtrAOy047Dd3/nMWZi7B3+cewhxvjtwDcycFZx5eMlw7AcOOEQgStuwQFYl4FcHh
KT0W9ivFGwvr7wn5I/Sy5E4vN4raP/3eIsFHiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Jh+1y0iEMYp5hJpjyM601CAcX5BlkwadDw/NxvoznQbqcU5lHaPt86IBU5Ow80VKBMvQ2pNav7xy
YiDJhNMDiS5LmkjPcKtIRTEpiRLEB5s24RgKTm2+lNEpDL9m/peqFb74+ftm7b0LP7Pc/3ZjkdI1
QZ9VKGVj+PyyfLWoVmg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OnGCO/OQDQa5iFBYV3b65BOVUit5SHoRhZw5mdP1Q6OYPwoZSnaiMaO/3EC3WqHZRM0sWEmfdPXu
XNbxSXd5bENCsS4QIvN7xNNShFN2+lo1Uhj7PIh4GXBPfNBOlVgug5XyzSoFefltXI1xw0CMLNmf
10plAEgakjXXdXVg6y0il0a2LWQSjAO3qFLu5GG7e71ZaCbQGz162OuTfIvmILI8wIIXE5ru3MfY
D6A6R16ImwPKdqDxyKCZAn+Eeh/q/DrOdFd3gbzdk0nD1x1y9adKQUQSQOvTVHD8UIKdGj7lOZ72
Rrov5ilWS878PL9NlWg5sUWDTWv2MQwFwaAkaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 141440)
`protect data_block
UelmESvAlWy6LgaDKEVDz9bgH1gULb5Ad9ptEWKbMuBzgqfGufXMBfMu/JsK1M/pDBqDtJSiS81s
ssIcQBfgZB3ThnAVVh9EEyXTlw+8u2p4X/xhoOxRbhQcTiQCjpxVxOpyy+VECkd2Tc5Hwf/UrgtU
7G/aTbu9YYQ9e9gqF1YTbx2bIIq1iHZ5V9kD7sv2vzBq/etNslbbnsWabbqnq4eYE3Bl28fW09nC
VuBeEoyAk/bL64lBzlcqCd9455ML5FT60Kvh4qWb3dQjHukiPBnv6kMWu7EE6SyVBRlbNAsLWKiR
+coj3ogoqpjqBYVQAG2a3PxuOPxFQWchAvaHM97nouTmhbzQzYo7sX7srZw0g35cyN310g3uG5ZX
4Pn6JOoYCcdlJSj5v8HZVYJHyFzMdGevmW7CRzP2NZ0ev/WaotdMZTjssj/aOvW5JwebrCobORD4
AQOPUKmY++u88RFVuPG1ROUuAoJ7wZwDrmolXFJd9El4wgge2VRHMlFH+4HEhd7CY0rFwx4DIlez
nRvMLBl/ksLaKtLi8Yv2pfgFIME9fDq9HolpNqm3nN926Gq1hPB4mQw+IvDUzHDE+hw5Tm+ljLHG
0whddbvT6iceFpTtdaTNpYv60pA0ZGfks2a5LYcR2eJXRK19QOrv47lnDfI5Bta0TykB8bZFe9dX
le48+JiA5r37KQJeFWGc5pbV5KgdaIH74d8+7WjbUOdkXOBVPebHyyym3GKefJ0sfnE2JJWom5lp
NIvNPdtqcpi6C6vV59OQeKbKsTnCCVTaZVKvekPD8QuK/fZCEfupVWRaCNRMx7QZ6DYVcGGGEkzf
tNlM4LzrTUfvElzUYkcIZ0vRBfo2VMHH3xMmi3qX7jpcEOgu2GQw2JP/VZkeZVTU88YWO1BejmFK
CInp1Llvfu349oQ5CNHHBAoc6PwcIcOe8mQy2jZ9t757kf0PlE6gKd7eRuEPK6QE+JuxtEi7NYQe
0OvJV3ucY3zcEI0GI1sERFw89ajB6Ji9JK+QC7aIXV+cfWJOxNwaWkpUYXoE+QASKSccZ4a2RHBD
mlV8L29igEmp56A+6F9SSr9JBbwegwKy6CrzTVFIQoTcdIZB32Iv9OBcTZN6OboN1FWexJmGgxgU
UgE9z79yZYks7M+B/l+zAcpM91TuJCZZngvNgZKY86teQ6xsg2p1wqVwGPYOzkX5R26JjktrTThs
thAyEX+7XkoeKxEJgqek4ZgZVDKpBrKojO1qjburCAGoQcdN2Gt15xDNsnrZaNI+z9jsekRhPc+g
lVUnwlpIsVKgQ5JMreRA19PbpFFNEei7utZ8LmiWo3BF2oh6O7iLAmQtDRhAXQu9XYQ2njj2McMU
5wVjbPimFa8b68jrLNrfg/gmL3UGGd0dSrMlagJgThdfHGtIEOVg5eAL5wDEcKPBBbb1G3dEUsWh
FFR5KK2MAhi/QEtNQ9MWn/zvB5VK13iKyFLDZeH1mbvRB6HrcQ6JTp18520NZ9C10Ow042o/uocb
cDN6nOkA5VxL1nLptjDGksaByxrrWu1dAtqzy/HdX3HDABQQgN6D7rZ4kEpElopnui02tr4v4OEt
f9/CMsIVQf4SsDaCcvsuRyi8upFSOx9WR87rbM+GI8DghPDJXG42oTaybSsdRMmZKpwsMT3cP3QF
x9D61ycDx/4v1yrRrycGjm9REj9vkbVmBDhcAWMKKvhob0jFinDovHu2DzBYJantwufRCG6sFBY5
7dEkH+iS0NCzlhUPKrfaQUc2UvLz4rTYdgBKbiriCEZufxgt2x22Y10DCpM0Hs6eejCe/TKa504v
WwbPTD/cWHqlgUN1odeuRBhSQ+Bc5iOsW/v3p0oR5v1NlyKUAJMeGIyoA+CsnVsoVFQB723BK0Xu
P/ocgH0fqhEW8RKnfI825sbiutOEz8vx8t7nmjF1g4DjKMTT6Ow3AF8RubFvP1feQareuplj18oq
2BaEH18kRpSr+MovIxuV/LwQWmOjtME6XdnKi7eg38eNwkHE4LuUYiVOfxD4Kgf7v+qVgQQl20mZ
xtKVvLUi8KaJl3HWaljcwIpuEAYc5ISCb+cyUZlI2lHJgQGElJ0TQ5/Y5KFC7DAAhaTJo6iszan+
NAlK0bX5KWVfKREk5s9M88ZuqPAENWmjH3tQxV2saErBlxcYRHFZeuCrqXgTTsxRUtIbXkYC0drw
RVGosRoVsgKXPuXkppc8JXndYEfZEeNu2KdRvYvb/zRdy8kRJL+Xqpdhps0xVAGM/baWEKKLDzhg
h+6l3I3+i7Tfg2rxd8m8J/RJMY/eCSEPNdbqBGprgUkOYw1Oh2+yxrfr0vKt84G8+B15QTWu3Waz
4K4f4suMqPLyYGEmOzp1OAlQvUWmQ46KP90/KtU9bFyJXTpVwKqFr9D4MFV+Rtpw/mKzijV+gY6R
GruN9Yn/xweWAaZcQU8U3Ro4uST3RPmPBp9nelChkIiofIeW3Huh82GxGKz5IrThi9jwMNrlVPkm
WKYj5eV1RnT4ODAt8v7wtDTb+dPa5AwbVJsDeuvKnHrRgq9V0Mc4ObYsQOAN2h1SeYC6vyx82XAn
QnEaiWmkFY7BOuzsxbcoKlqMq9VCl0NL+pcULNGZe1R2UbNmnnuu7189xGHiCfjeDbUQrDITprWg
2hfIYI+fsCqJLnhK5CBWGe380AJNhe1A2Pc9TuNMb7qXUvifimV3wJNcQgIIPXFXR9f/NecXGnNc
exQExztgWyPoUTyUfPQSb+zYbQYnuO/GjlmHfzgNQZtulnUrfA360r5sNu7z9koKiYH5NVKMkEN9
2Wf5gQvK4hdnysH0CtDCMJQjukkrRcDvDU8I78WazVliMhWyvwzdJOt5sYcU8sYraS45EL9tzk6T
FDQpqv/y81J0sujZl1XMYmDGBEgzTZuN/YFHuYgwCCqveOVGwjGwk1XkZ/dPHdHp3AQTetAYUgbX
F2XIp8AqkgWrgVMgyqV7nCtwhliyVLcAp33UnV9NJAKe8Ri3aVTXVavOMX3jirfgIBVkPbKRKoeY
OAl5d3W+NF6wI5NyZBr4hiUmy0PY7kBZtiSvDJPBObZLJ3EQgnNzHxlDiCpK4DqYDpWG8p3w5IEq
hS2w8nGM/rEhq5ltYP+yZqsot9/gMPsRH40kvW0gBeZnijDN35xr+ZgKeu7NLFJc7q3AQqz0HD3i
TYCYNfpOi+5+sPnTWHHy4N39dUttEPfqzxrWaCadhRB18HicY8HdPiNMYx7xJzXqrX03ioqD8Ro6
smcohSNuT16YIUPZQS76TlEKWeQJQW1XZ6GHImhXJwhHrkOcNs83noGIH7JQb5ZcemhPem+QERcS
ISp4s8p8a8X1EXIbiVS2bK2c+DZ9hiHiq1/T9G0OsIORQzzrc74FIMDN9WtdvDNKQvJGg4EtaoDp
gwZgszyi+XfsCw5HT8fPK4txoVJwBCrI15voPSg8xp4I49jAyvKsBqwCgdoh6Pdtat7McqWhjL3d
b3P5aBa7U04d7ZjoE5zDLkLzL9k+1NE6b5j0IUiTJ7TQ+psemeixk/PshZd2+s6iLb5Pu+O5q+R/
PdktosjNUPy6BW0Ycjjhy7+ksMV/XGVXymM7E4GCu/Nd5IhbjXEyv6Mu52bB3xOLBpOJ114TBKBN
0lf+lVZBEFLqRZwTezVMjgh9O6uSZVEwTr73SKhXt8w3g7M4cegHQyS4CAQKczA2ZlfRsQ44ZkQe
q8tjHVE/tbcQKLwDLlJTd4KL9nC4mvL7/dk476OOwWc+fnxKiSs+nsFNXfLXpjE8xfTHFI7hrk38
IKUFIe4nSQwEII+4RKXPzLrsKK48+swPlrP5rY/r7QmWHgUbimd1HFnwgJ3Hff+JlWhzO7JDhumi
cPlTjJjbO6BzGmUsaqPHNRwHLZANLsv9FdupOFBWx7Vp1ZyFvVCJixxdpg59eSoY/hSvDtbJpbBq
ASBczYqNnoM45ZGqWNFh1rZ/Qk8nwKdmbBfN7zE3mXdiD9YSqm1keWe2XUho0ldzHyweVxos9Ser
Z25VIx3eoo+GOToDMy1O3c05eOI1f/bobVbEfZaOqMvpBq+FhKi5RM0cNW99cf8fH2XPK5ch5Qby
4nJZxdyDAun/DpT+aC10gyjKA0JPxeVk/eMTjcgv053MzvMQIUk3qO8IJF0QqEFybnsEWJJbN5BK
hXNLJZFImReYQnWqxDCKMxouHXAcV7KbV4ICdIEY0x/X2IFdo/L8EJkC/h2ffmYORLVPRSxaX7Ng
r7C3AKfs1lS+HKgbzGHdUstbLU7ovGIpMQrM0pOrbH/e9xkiv4Bb78SZqr9SnKqo2FMTrl7ay84P
y0MLgrysMWggFZdovN7CJxyn8Ac49Y3RMgi9T8NML5eOD3VClA1fUGqZa8qhbbeXO1PQSIqPezAn
utbJoS8uDuE9z30Mbocerhy06CKAS7e9obXapRcUcAvRLeiq6QJEIvU8f6jn/s09ZWnilAwfw71l
FS9aYF5O3g5ouLawphA6XgeAH+kl7NMgogSSwk9POlevd4hJbl6FppV/EY/er7UTUWGXhMUxkuLd
cGqUjTyc+nUeJkD1fW2yF5Be8PuN2qURoazeJ0Kj+otfIYLU0MW8WZF2WelNgYt7atoSTM/ZJ4KR
40yc802DeGSpegvS7Kdt4g+mRJK4LvdVpLgg8yxihSmSLN3QjA/TyuIRthRQEKeGzer8L5v4w1PZ
Y8dzKtErjSKFSoNAmwqnwYzXDLQZzxjT8f+IpS4yLeJUIwvyIK6GOUJTJumigGu9roUp4MDvePU0
5flf/4xatR0ZByr/1cYclde9tgyW0iGKXOdvIUxGTkRrfCtjFNjTKko8hCLJAfFipNbmAAy/fau/
nWgFVGaj6Qh5GkiqMY9orEIBmeiDNTdWk4Rhu3ov+rGds/WsXE/OVnYV4tktyFr3SQeLAkciDVSj
CfN4p0XBfV16zYEs0IRLEeEq5aoXpqDF8Es0r5ilepQUbtnJ9fIvxW6G8qMHqizcI116iLGYm8rR
r4wxFYionNCmIERMIw9h3xFrEuc7K3HURJ9kmAqe5xtpfErJQSWrAdHgy6FEUDmfOwOzQBLpprAt
O+p2CnqFQe3IASBev186qy0DNTR9/THMIR0T/CmDQtRsRdkmeQqwUZJujDZLMzHgC+Is3zgUcqvt
F+hLwa0C1jsqm2NoZ/BFZxd2CrYRgCQvhnnNcKkbC+UMClPJBLjX0HSFYoQygKq1/fpWsMBfQwCG
VwBQynB7zaMRCUIuk22Nbpx2VMlxfbXulnsQuWqMpZp45oRLT0eE2uKmnNm6jtmijPrwCChLPwSL
j42sKt5W3b5ukqEdpFd23YOM2weDwwwTo4hol1nAuLi2brdVku0/s8IVUUViXNdInWy0Of9atO/l
crhuykk9m/tnrkPhNOlyS+KpsBPVKPJCIzuGNsI86VCU1ewSYYa7IFfnxA0RgnkNRIGQGwvDgXqH
FaXHnbSa15I4PAHic/tTJR8mudZlJl/9XnXRtgEK7i2uoTKomxkDb4Yz4L5jUIcZWcZ1ZKAlTtRx
ybldLP01PS88tZfYS9NbtxN/D5C8bC1wwzuWne8H1ttiiAK8nv9nn8VHKTRo4xAxcV6KjMuDD3XB
2RT1QTdjDtxwRduh8EMImEJPC4AtmGSbcyfdx51T82oBmc+uQFtFPpv6xEZmt2Y4OqbNvR/S+v78
46uRxNzv4nUHoBT1F0SURJKhnR1P2iKch0lC4IHGjsBXFAYJaDz0yUHMD0GqMHWnsTwGezdP43Of
beiCa/aQ0S1NkMq2Yb+WGoEravNrHcNqdGgWGTfiE2I5p+mFc4NTHRV0qZkkw15dTxL16+ugXAN3
UrOEZKV6jKmMgtvlF55KSK9lE/Z8wSYrZJleJ9j1QYEmqJjSgtwEGtzH38Hwv6MjSwGeoyHOYn4j
h4N8mn3mQs/D5qbfXYZ2hnwZ3Q2g6qPWU7cyx8fYX2r2tQ9fQ8L6RnHoFti68M7g2vHBGSkuko+y
WGYeYRI85sDKRFbZMQ/u859j7aZ0gehgo0fmO9AHZpV2lLDI9zAgId9E9OL7i43c6E6wGZrGr+LA
A3NftSYKWlAiRneqg+E1ktGDKBYdawd0V49ziwE1Wi/xDQ9H4eENuyBi6ZPuUVL35/cGv9nCw9VM
RTfiIY6Ta/XmaNGLbk860XSNePhcMjr0pE5ECk+JjQjd7cR2zhslM67IoLDE7J/MuEM8d0pq1lY5
StSlno4DyHLIWv53iQJ32+n2O9ZIaN0S4EMg02iLjUoV+3BYYFPAd9TA03BBW4aKGkMP0HJMhppG
LyVLnVsD8XssTfe7LwbXMPYc4Gb1hBFN5V7AmjZORfmkxKhTEyJWMuokmPg4RpLCSFSM2OTR0Pm/
xYiwUCuaVSlaOi2jUR0IPoc1QBJGpZQh01P8R1HoeQUxmgivdxENWVZoIgTuLeKkcgZLl2bh3ju8
fEigek2Vtmf/k2NF3mQLe6Uel6WEY2r6Maz1Oc4Nb6u29UTDtE9NS02d4TOF/jacdYaq6J4Mb+NV
vzBJekcvssh5vv/aYEKIsUgJScEwJ0JLSL04Z4RwiCW8hNwYN5XaZdrUtUnWt1upbrnmrzyputRi
tjDTG2VNINzbJw2dnRx/OY2hJQ5djYhhTQakWIE+nMl/66L4pMJV8++AXsYir3p+v+/e0rLRrjpQ
8xwdEK3b9fNQ0fq6Ig3Co6wFPwimLCcOexn7L7BQf3labVb9QnjsWBz09cMK1Rn3I1JW2W0aiimD
tw0IvQCQQQyALDtagWlw7hXD+rNufjmNWG4uZFQNpLLstPfzb4sHpDkDbjJGNHsRFVwTXIpNPllI
SgBcvd9EQr0W/UDa+qPTDtyI6QlUanjM/R8unifuamDel0ZDl9SP998BnCEiEmft67hXSFltCtFX
ZTmVobEGSdeekLvyBXTLAe51PbMcrYnTREnlGHlH0I/y8gjRDpt/LORJudjITqEJXSKEGuFvH/ez
fXRCAxaBdVWmjsY0jFRb+NscvTCHkGc1l1d7KakwVcNs84l9ezuT4j1Z1IDWaXBdDQrKxyN3gf/6
3sT8nBn6Bs6MsCfPwOvkBuBMkZ0HIMPPJWHAkrcbR4dljbzXkqU3Qifdq/+cp6TkTeYVrqCHkKYo
8IuIHCpbu4fpi4EtozybjNbMw2r9yJY1sbI7gEdNEQkPd2GgFdU/JJ6WfhLolZMAY+XJ6+NN12gr
f1jLX03TZBnM5QyQe2DBDW/4uhCtWuMj0yhaq8stxniy2kAj4CdkbilHdxJBWZss+wxNZMNVaF+u
hh6ZudbDVGZHErwGy23+Q/aE7BUbzzeZZc1uNs3FNDPezr1DquZkJUyJA9e2BYGiA+hTv1bAV85h
GqDNuXD5Ohh+qcu7hKRlcgUxOU5LEq3R/pP7nOkfliABerMLD4GVrhn2zbQ/0z1ycP5Mh4PFdGSP
8tZGU095n/SsYrxQuJUBQTqC1FuXVPU6nbDfgLQKOwslLERQq599oYIDtPchMhpJZ8zk3ZmHklSO
xBuc+FadFhgFf/QGMqWKWtsLMts6kLRL0h9LzuxIeFWwt29tY3r6Q7b5g14BbW0aM9YWfkt19Exj
SW/1fXb0nZp11qx2g1dW1av908NkyoWnDM1grlkx9PaSjDeH/l2pNwNgAzPb0MgOSXYbKLDOfPK+
slYNm7FuHDvmKufuWXmbIlZiuP8XMsRkbK4I5i09STXRq2jTeArxSbglxjjdKZlwOeBrXooCzdXe
lMk1nilacYc9U70pVhP6KRn4IFedGvem6ZdbIJ/w2v8fdg//ppCgw62oRm064McnHTu5aewDWBpA
mHqwub99zqDjX45VPe/z7be07mjSBCwsPTSnxMuw9xSlGcvUNTho32+ZNwE7P3VthB+3frxNgWdP
BTw2zbS7jcy/ZNqOX7YAfqDP/iME5WG958uhHG/Vu2pQr+YUHB4K2upI+wUrfC847B4ek7bMJo8p
36Ur9MLSxZr5D8KpKKxC4ULKGnOthRMq3zQXY3QMg6RYIw9UNib8QeI+U8aCk3+8Oix7vQmtRS9d
/Uw+5YcJjUkgFVEICwIFkqvnYH/QKt2eyUspjfFiRtNdbXIxoEos9LU50LM7GVZXShUyKeczx44n
3alC9rx4ueo8Y+m1/d+6BRCgFmDBDnSAxrAhp44GUyrVoWb0ir6rbvPPXfs5zoNPy+Q9Yt7GAl+K
uZZxkKSiP9bNbgUmvWiSAvpQF6lq7MbVr8ClAw6+HEYZ+d4a/+RwS86w0aCf2FRnY2UM+4Yj8C/Q
biMWVMzEQy+oj4W3g299BpHmjOphPy6MGf97dyd4kLGmltBpJtNDAU7hzywjRCUor/974g6NgJG7
NKqp57nTf1iUzqVY+BDqh3XzWLBlq/QKX96Fdqh8LvgyMUMdbaBtdqX0gpQ77x4/kTcB8SOJp4r/
FkbJDe2vTD0xLi1tneomnM1EZhF7g9PJ8qbm/nGxsAXtAr4gLv81AE5FX2J+jKMqk7A2+OJYSYjz
+0+0z0cGwMuXq1xk4/zyVh3X4l2kIvUy3g11Tl1upm5iKB/iBM+wHruyMf+9Ib0y43ls5hm7TLHw
LeYGUwc2J9HdPegNxmCTIJF482uuOoftD9MKv2fjb7Njb3/Ut20JoTFRduUbYFQ+uCwLfpAVC4Sl
KyTdlEMeKLH7gwJy+3QYI22hODpcRpu+TG71SBrOWOA6KJdjpVC8beaXAM82LQAlOoSvz+OPlArQ
E6mkYhdOZ4Fggkfj5NkNwxTevqZ8jeFVznvsHHd4y7GF9K+0zKc/5h/ldX+6qsmr+kkImBu+6Qox
0YPXH7XYFYQdFCF2AjasPoVwpzexaVEQ92base+UHciGc6xf7qUGbJ1MAn6NEu1kKV+V5RwmmqxT
5BbyFVBVw+DhC9B7J2hnOUJyXFfK0jzdw2Rj3tydKOC1f/92yqAA0MuglwagWJdfimpjg5rcHB1I
OdX47oSFgkrdMmbOeuNsLiTiNqvEDpJNW1BpKv6sOLSCRqwLq5xuTKdxEAAHnw9p0gFkd0+E9Ewf
jdat9hBFk7BPPz+OJAL/ApVVbFwaL0AvguVYit945+wL15x1P5U1nVngxJfbhV7UMx+al0zRcDUs
a4dCl2iED7sbDee8FWjnNtD3Y1M0ZES51v/f7DmxlUF7ItG1nn7PYEKeT7nQ8lZMncjp1EHaY8Lq
6mldAhOr/LEJARuMrYsernnSu+28OSWnbiOpHw9ta0iK1fb1PlyoNsKvtrcpDOpaen1JGfszplOf
Ps1N/fyFquOtcW3aSGvFaE27ZJOVaqARVH13N9pTjoLhadEsqXRonPQAG+sdK3ZjdBFDJRo6Uo9C
vhFFK0/6JKTSbx9NFaMqSYIQYFiD2vqtLfqvK1MLvgsdForC+L7OaVKiq92tWPDVmfKQ3ECLJpjv
NP9MwEQgJ9UHKkqnqK5HpqyKAMY3omabeJ8/JhOwM2nQTnyDHONyqHaT5X7eWiFuKX30YjdJro+B
c5P2fj+8ljeRXUBnn5bq1f8a2g6SNrVo+vXuRGNWfZNu5c+6eokiiorCarsg/BQJnlM2GlA6DmlF
cg2dJvklSNylIBsVRUCobfFv7SYJEXB+v1dD5dz7fd6amj7xtciI95sNMTa+EYpUFbnYY7Rke1Pf
cA/7dUBzCyD4vfPnr9SHKvMwLxgAFJkAYVvo+xaqVIuUgQog/XZdtpJgUcRUG/RGVnTSy2Wl3as/
0hlamU2hXC5SJRy9EEZ6kYGDc9McVoEdhho7Q59qWbnFs/vQI+HcfZD8opHD5ffnLNVN5ngrRKYA
8+EMaZ9tKEwQTdA0Ne/cmRwVZdQKNr85y8L/8UCnbkM88n5gM40SD7wTJhm23+FnP+YiLdP7Th/L
iOfYL6Fy69JC28uSt9LpT8CzrX1IWeSNhWKDNbHuUyIgeKBPNDAtZYBoDbQ2nQrVnP8Ot3ZqSK99
8vzSQ0Fb5QX/qclomw4Vvllg7EwYScwFliQNEuvNG4/saOTfc5SzzDdHx6xJpy59acyb+LTSvC//
cZKRF+aDFArZw749uSUEMtTmuYwIMDMPiNqxt18gXpChk5157LCuj/I3zEkuILXKpBdhbl4Rvuzz
4OzjVaxYt11DeP2mu11uHlbq2mV/Kmwk7Y556pln4hkUHn/Sk/cBgZLfrBoL/kz2vmPWwYADwxG/
yFywdUiZuHC+Srajf04hWufpPD26586T47VSSeSkMKeSOUzEAI3nNzp6qVId+5Yjvy4h+NHBCVJh
FfnPz/alP0WkhfxTK2pkhPcRTC/XPiQGJftFhp6kb8XWenvTr/tikKAu8qskJa9aBYFAZxs3Tqrc
wWjFMitLhqB+CjY0Qbiu5DeqPDcHfdmf2M6L1dOWInHbyCZX1aH/v5MUtB3Dl581hiN889TyEpbe
XM7zpsklFX0tRnotNC6qdHJLdHGSUvYwJLE2YmDftdh5tOxDlw6nKziFzM/JaLnFmt+sNY9+9wYJ
B99VCqONw0RsZG3oi1Nmhg+bhPg1QJ6AAaXY6pfIrIaP21IbY204hEP6HypxG147TkRz93mpiW0B
6y0IHQ6Aif+zoZLtTGyFkYmA6Ncis578nCsTBKxfO8fw8trGpxqhEBGhdUnMymAbcBhGgqFAYdsW
A82iKSClZWNveqx1s9f1GPVJfzy20d678HpLh/cpj2TeiaivpF3V92S3Zqn9LkFo0VCOtxgxU72y
V2XehouZ0p86R0Eh9hlYk8zAGAkL0LEDP2Qk1GCZPKbzM5rzuNEiKIfv7WYncBKQFsx+FSxKiDfK
mr9X44za02ByiC+LaGAe/+0nl92H6R4gii4vIN4nO/VIV48wBw0MGJ4BQKJh2SU60fzoTgsbpOp4
6TxpXuaYoA86j5HU2INYOYLAYXc0PnS8ptW9SGzzhOSkLrWRGjwIxnZES/UCEL4/LWe3TytgJ0gj
NgDfOHtTp04bCM+gQW2T9dOv64F1Z06lGl7uVpLV4t2ivjnAHdPJ0ld6fPRfGBbTMM1c9d6ZlkNz
ogpvF+sBjb50HUJNE0xJdLIcyS4i2MLN5MNjiX5UMcAYUx3uVK484w8ljdTDMeQQb9+cVs8ZcXqw
wRY7R3Uwfp5GeVRE4ukhQlEE9XebdUNDMsQDonrs+aB8nhxVWQ11cb7jD8NM07GNSeqXv/OjMTmU
P0yLLWAy0WqLlTt0X2YJ+QIt7GHjOsbhzraKFJlaLuifk5av3rZ+Iv0DlyQ1UbcVLkNg+V/vcOaE
iwaGG5l3V9DRfiEnnCRob1h6GkioaT7wAawkzaFxpP6VfyBeGIt3p+z8vyDfrTR3tNeL2ChXcMrV
l930a8if/rgdHpcV09WdORBm9VGY9PvENXt1zTCx8YqI+yC0oQTem5vJGts/cnDrV7OveMsK+IhP
aOavwIGJC3KwI3JK7iZ78OPrKFCraVn1FSpuJGztBdLvRNZrXyoVjVYMzh3RX7uFNPuWCCZrNU2P
W2Z0fgBoL8fZhzeAB8y3/+jnwzhkBsYq4Re66+wgFSIq0bzybt0v2wPpSNSezF5OuAeD02cJyxA3
rNhcsi95WOtcrkhDjn31oib2OtesZku2CDGdt5lrolHOsEx06pkGZaChusJYPlp5oGP+pvwGWW3O
GXINg0DyokdnEtTPZD+4YBSzMAGBwK1n1fLkrkROSas3cDkgag5YvnwBoiLx/CxFfcA7HSWOppxI
+cXmO8PWrRxf1A+h1VY0Hd++CvK2BYQevR1eoGtzqxsIFJop0alLkvyqNdgwJ+7keSdj4o2nsk+J
MCDxHoaaNUr+FCKzaeySihOedBK0pIVY4RZmd2I2Ce474y9l3S9a/tNH9J3GSZd1Aqwg0eHIqQGY
YdR47TkqlXwXuWgQu3fAx/Dn+26SAXumGSJQCBkvYX9xqCTpcN8dIG3rKQAyniavs2Dphhbk9FD5
eLQRo9HdHy5iGKBiN/ncr0SoxKQnvEkzW8uSE8HGSkl5msj1/w0w/B+6Vcd+k0J7xSgwugaN6R5Y
eGJ8aR+4OqV/ptc/XASXKkYFSuCSbWSjEwiGxxhTS43cr3wAy6oB0OQB1Mrmknu1fFH+fpQUJUZX
C9DcXBO/EWv+BArB/CdwmI+ByJwkU8gJtbBXH6UWsV/bGiqIaqZK8dRX+hJkEfo/kcBBIQ+6egjE
AAPSHmMsoJceC3wlnFm8IzZ1HtPuYzzQYPHtMVjnPRD1qXP7MPVmSVmoqPI5RRhoO4lur32HdKa6
2MvXR2uOc+d0GYujkMf18BnydNN3RaoE1JzBur2LA0JOIESD54sggcioV0XBpLqbcOpCam+3uTV/
SDbSr818r6o2f30Ww8VPviK5CsvunxboGCEMTPU35UfYLUbxD87svpVpl0kSjvsrSskVcGFY1sDK
xRftUOYGURxMY0SP2fNI5wKFuhoWDvETgbQvxpaqyukJvf7aaWL9EhpG4rUO2rToMT7PZZq7/DaI
ctxzqH6dK4UryhNjCcLkvjA53LltoTF62INY0wsXF+fsJu3E95ENt+tT5wmh1Yn0YJFKoeiBhc8I
oInaNT1yORqc40cTNf8Ix+tfkLlv3FfvMt6IaucbCAobLlkuTtu77tiQKFYULtZhczF59VdmnNaa
lo/QXOikPXQj17uubyd83oVsq8cLKKsC1OGiXxuya1tQ/HnKwAO8AeQ5aAv1yrYiYknao6Z1DsbX
aMGPjg+r56SNmDs3ez2aL5IXGAv+W+uTfP90c4YozZW5izQgfjkPiykg+fug7tdk3+djXNRwdN0o
LwaUS369+OrnY98KIFZ5m4muHUwvKzohs7LeaTaG1OXFRC7pPnOAqaqTXQbcR11iKQi2OZZDN3zQ
tgsZ1mc9pco0EWo/XnQjpB5rH6AOnQJQ6azpxErCXBpJEE8kpIRCbDRYjMBY9JoFAliTAZ1Ce7Kr
PeNAPpJw9L5Kg6GSrO8AXAYRHfSjZaM+yoA9yJlcvEJh8ax9HzRAKYFtB4etsJj2KbXZYLIwGBUS
p3KN/qBt7hGx4zPXxnRt4APOX0r0CpNX+rnarjViPvdQYEO0HWKhWZpLNb+wB1cNL6gv3EvtVxSa
JPN00vX9phAjJW9/gPGo7OXjCzq9ck9swN9gB6mdVS9ikC4d8emzL7v4fZWN7O0Hfg64bvLAFRT2
yp3dRFZ/u6/fnFZJwOx81AWEgrt1LIij3MTc7VmdfsQqMdRloGlU6C2Ux/EH+L6svCDxhi/ZuZcV
OsB/BjZdzlZ4Z5+pZ7b1bby1UdVYbottPiJxbSjGLnyJMjlchVPVvNQM9pjDXfOb1QmLtsMhIzg2
bcHr+XvLfLHHwRqEha0qZJLWGG0G8LvzU8i9o8dhgFf41nPsKfg9xZk1dTl65RudxvKBLyL6GYmm
L4Ibqc4gQV4ueMutukkh3g5AuALX+2vfffWnPzwC8QlBAlkz0HRMiUw3crhCgBIw1AMoXPbcvfnX
S+3UPE06VfCoAkVKTEIc33heq6Bc81ljDAXrJbULcp8VJ3MT7VqARLbs5x3Z0GfJuATYETtAJDl1
3P8jqHWesnWTjqYLH7YhjnnEdw92OPjV1RyrXsfrwx8GDTxZIt5WNGSDS7ox5Wu5iiq7cfok5raW
P/YS3l+LyIc+G1S4ys+f7Yo/c6tuTe6yhfl+kS8Hhv2a+snEEpvIhS/Dhxup02cm7zaVkTt06B00
l7uE3kRfXUAF0dPkHXN7KWbTdQtEh3XykUszz5xF7+oWTZflQbTyDPYDQEzCi3xs+Zd8ONSkszXd
684v8b7q+wnaQEtCa9ZwhtBXTbHyuHQIY4sH74qTcKI2OvF4WV5P2I6hX0CostsFNsPsdtJDF4I7
XNvr5z4fLEOrLGAm2Ss+STOPzSu0s8ujfvIkotRdH4mY7Z+H8hhsLKtfVBD6DfQL/jIurJ3k1b/x
VcehzEoOS9Tbljw0vh79GBGeLtIMor86W2aWo4urxNq5ZZLfP1DolBRvkSAo2vS6yk5w0MNAjQYa
KoRgxjgO0o5pdPv2PnrRcJkUb3+fUTmaSSrbCxcr1EPmfVoCnbDCfN/AhzAFJq19uuPJ3zEDU/b2
2YMNupmWdKv11Ua8xYbV+Em0ZflRQb/+eiFDppWxIdu93TPOmpHpeVD2+f5NKmbc5qLikUTqLnZ9
hR9GGsUOkNNfnGY3o3ATOZi4vsAKySj0GtEXEQUQGromtXCaioU70zLyjg6H4uNZ4O3E902Cdmvo
StNDLKD2DYiA5/R/icjPI5T1y48ERYkF9qzIgFqrSZ6LgI9SFWSlBlcgPJU2rlQqKnvkwL3Cbdn8
iHLa2unegKWuA4whWwyLG+4TmWmydYpDCshAdGDrxIWy9R84eB8UJMnru4BYSOwl6TFzVOgrUyYD
CMCnKDm50X4OZfm4kI88R0GborIXB7hCCfYPA4DXiS2SwZbwFnGrNmbmlvRUDTdDKm78MNMD4FRn
x+5yv01RXLDNEtwlVqFzULK+dtOQaH5bOH6MNpbQWygkle1kRnHg0Yy2PBlb4dwid4FgFCEEWQmq
xg14a/qiCNF1jMNv4B9Kthr3O/FsEy1CMjVLVQHuytmgI4s1bHa9KWqK+t8A9luqB68dOsdwUz5i
Uqb4wiWDmsmLsc/VV7edpfgKUwH0LIGKiCeZN1JioFI5bqcZPv3EBXFoElzNUOr/cq8rFsbdG4aw
ZbF+j+cOIEes/aLGV0ExEowePp0rqxwgeLMcp1Qu1jadeZiJcFJWi9axbDyMcWjkEvaSbGAjhqqW
tz8zvCV1Gkqxwnb556+Rb8+aD8fpvNITmVvF4nttAL8PVGPnIifS0x4EnZgP9Y88bh7lOzilJA3H
IUurFf7GlgjyrOVXq4hQm9PRAjk/ZCN/SFRDmdMyPWz23Z4bqSuVqTRuqRgVDUMxTKyWEU3UfWBZ
hJPB38+cvjKVUKaB7Gmq4KORCqHg0CFX0mME7d3t2A+7vfQ2USliD+biCWRdJEyTKQ5uZbOwOAkA
Tknnmzb+BWfJLIQehddU0U8qKtbF+qunxElw/f524YBoVam7xSYWkk2bofpIDGRwNkI63qZlxV37
dTdHEBpnOhNjb5urw5PL3NIArFjS9PmpFGuOXFbkCPvZnfyuWTwJNVZ6sj5stj8ozRIfkYAsj7DS
Z2LBZfnz00RM4VzshC1hZbR0oV8Hrgj1C7bBfPOwrhKVs9R7E2u55vVpLzTwSUPWj3v0SNNCSZPe
2eTehCo0MUAtdj34iueml50mhz705kCXNI4A6ynPYq6bZe7fcbUZiVsvgPTeBsfpmCYQhW26jCyV
8SYnD7oBmtVQoVju+Jjd6GzyZlojEArK0X9NTpLyoO1cFbHXOb80MME1Ob8Pp/4xiR4GnKpqMXm+
KNHbY6Myejyoww7co8IfvUZx/uIIU08s74EyMzH+L7jnvx0Yr2m0diy4sophzFr0W3kUtZ/Nho59
t019xnLrE4JjHislI1O0asjbybJITxN+uTfyKSwdYrGesPLe6CeRyjj1zQJ9HmfDZUAschrOUf7T
Uvi3TKlkPL3fYVAdtzh8+mPzYZLM3C9iV8rHbxknHMzSdC5VKLjlhvUqsJy7BJSOXXUsSzlUSCOQ
ZiNIeni9FlbGmqZ1JGqXBwXkONcVI6nM0CTuoeto887su8hdINZif+XpQHMt6rVgyg2HFi6op7Q9
hfCAyKPSpWpeJd2s+fTn9wa7kiRiK5O5goaHwzAJ9DC9lCuQ3hu24THhjSnitYheIIzzLI0YDmvI
nnuJGF2ATOtZe9VzSTavSxGifXvztMXuL23823kc2UyhOE1djzYOtELLm4XWNJdXpV7ToBSqKfus
Cyg7GwoByBHRPJOpg6boekAhNKCXDS1A9aFh0dfQyD3P/sX/jVypHkm5uXFlpoc9MGhowL0brg3G
wFd8feYdvVRFeFzKX+GmB3jNxfMsMiQl7wlL5/DdgE35f7rlgFOSYVXx+kudP6OmftMr6lIO4NVh
nnWntML3D7k9vGqKpUhMr41mRjH4ldMU66WehHekU9bSEzbRJhp5disHFErgIFmfwvdcVQorRKWt
TDIoLmPJyITJWPyJDvW7w29ZiMllzIgAKfvKRWZ9U9RgtZMivtOefwcSPYsnqgcfyUBtOngLMIAr
+PdVHKS82fRyo+nMt5G0zjOv5KveKwsHedpuDhLAtIUkrJyL2pl/7AE9GxrYywuDyAkbsMVEoZRD
XPjF5C/A7tcwpg/gR6+iStRPLOENRk4BuhCYZHGW/DF4LnkhCr7Glf6dmEULZPV3Gqp6m/B55d4I
KnEMR5K6pQKPsLzyhUkwQNCTqMAe7yX7MtM45SDemLfDLzpn89DrSGfl86tdInRoReTJ/vVPMzvv
nmlLS84NjXxfd+41b2QPK0uFhgya0CBWYCT4aephTc69p0f8bsP8D1bw4e7FJyiYLBSMlHlMJ19y
ll8sVwbUR/u3FFv7E7nEhpIDzxQE3e0nvLwLVVQtKc33K9OEN0zn40sOrG0V1FFeZA4rkRcxqBR5
9ZCoScPsVrJtrSHVCr1AfWzaYZ1esHCkXsn8PUmZ1hci2nC3jBSQYoc6LZLjD20wRVkRgtf4CnqQ
2+5wHiYCpDxdasE17GHL2CT+IBBKkY6Uj+B+rnmzSyGbgF77hx4N+i1yvkLIzL3T+w+wfnbqJmYs
OdiE7GjLD9wF3WIR+rsz+ZByau6Rvvta5FW2hFN1stGAougOu2AA+dVAOOjwdEDihRsV+ZV2q20D
8mA883jBrEUcy+VNLTsy/fm/LRL5t//sofHO8186Jy6ffx9VC8VmDu3Wll6lpO792F8iGNvaHxSA
ihbKaTbgbhvMp2TZJ4XDm7dYmfTTFOjx7BLZ+Uc+6Rf395K92fOuFdqlwbyHgogeM2bXKLQifJpq
ycoCrFDvuGsjbGtu3CxU1eJudA6rJeK6yjyUe8Rwx1ZLKxKyru2nKKHV7LSFVAFwELdqALjPNx/5
Z9sTggeKwJekWOn5iRUd+os8xeBZWVCXuHs3k0lsghavoT+Pd0g6vKxlI4vmjZNm0lmjJ0F1xGoj
577Ba6PilfMnauW3SmmlO19BdzebtS3Io+4TvH4XejGm3rbYI55tdCoMGCogW/WEUCdynup8kpAF
d7JAWlX5bGT9ni6WQdZ4apyLCqXysT4AF7T5VoR13LJFS9bO5OYvGTm6i72HaYHmehvc1JrWPNFV
Cm6FH0236wTYDj9oPAbgmicAIKWQbFUOiN+DYWz1AszVLTia0Xw/LDKklMNzLFPxm3y55z10Ei9t
JtPV6EqVwxDtMTVSRirBbxvzWHs7tgO4/Gxv4llrK3Em/KPtsgGOYkMvXATYjyl0KwHONNn+1S9l
NbKFPXBcMNHRtsVToqk94VelvjLdlFHBgKQCVS8zJ9KaV2GUlx/WDyT8HsKVvfAk+RP2wmImMCgr
JoK6P21BAjlEnAXjGrR5HU6Faq3zyyA8W4qxcBn9aBf/56yKGvIOBRKJG4FH11zREd8fFCiLm17Z
KCs4Zk/JzfHOyZ+FCQ8jK2snfH2PUMuI2RlV81RGQMWK2PX/zqkJJHrsJD5j33FKJdz7UE4jLUV/
8uKj72epGO2dbp2KtA2qTE5iyk0VMkWXr/cHopQgGqkznOYZ33+WugFBvjdLxbnS9ugHPye6QKon
HNvEZenXZWZeCbmE1TYLf9kKE2r8EhhjB3CxBQ0GYHEEmDEdgYbYzTazxsZr24joIqBSloAnzH6E
Nto+/VOJCtUT1gPjGRAp/3/iC0eQ8BD7kNXJD4j3I0mD6vdTGCPO9OTQW0SSvMxUBGN8oMFCgR9Q
PFAxJaIURJeI9F/hsDca0C6Vofdkq1yobH4xeYq2yuLffjFW9IazzMxxvUMfJeJ+VT3vrq8GXyOY
ndTOSc2V/cm9QkS6DqTvIQhWUY/LHos7v/I7cfgzo0Wi192j+KPYab+eKZj/8jk5ZzGYDUSqC0ir
K8IIw56bsQ/itvfC7Jk6RgxBt+VhhbKyZ99QCqWvH66i2TuK1PWNPKfZIPAeeKIJKNfsnQuZfcAA
0NOUgrv5HVOyM/UO4hs+RhOMtd01meIPPZ97EdJRilPV21PjfjIliaxteNOPxNQSSsFiGF5xq8uW
FgAowYhR3rTWM1Io7+vkt7cQ497i0uVB9IjOqMcrgTqvcIhNoqFiFRN2IaUWucUeuSz+wwpQeS7a
UB06m2TV8f0P74ioBaP0PTwDJOfWFcV59XRQZ+ykw9ATN82c4SeT6slXpKrViLy4X+l8VFFlbPPi
wfb6dV1pghitM4zqv0xB2O5uevkZ97/wRyQI3+3LbwHmuUhFFwEUK9oWUURFsylT3UgtuAmJnpFQ
IWQgPkhFHSM4r4InFD5n63MAbpsOrCeKOagd2kSI+7i3/ByuO+zVveEigBHv/YQTCq9izCuRBUET
Z5T2FZ1zdgtBPJ50JmmCUpDpChzNMAsonCzoi3r2fpcumzE4pTbMR9LTydkvq2cmIfoaOOYhccsH
I3DjJtqVHSdThbFjbGDqcFVJkw/TFXPuzL17V1FebLU78nt63ZpGCseqcLBabWWzi0CVSJ6nHyGg
txhHl1XX0Md1vUjsn54oEFGO5EqA93K6MFyH1+S2vPa/7T1hUyduBmFxlPahV2qFoEyeYY2QDH3b
WkLy6ZkuV+JTrmPfobqWUClLY+mo4u1NwrwVPiBu/3p/1mJYus94h39KCnMxO/DghvDLbKL9tYN8
lhIwgtI1xnpl/E3DL1h7yVLeBOstMw9vK1p/5OktHH/o5Wf02hmhLg5vMLe52AxjyAlxjWWNaZ0j
CP+RFGYdwO7l/Uu5gDgX0TXE1Kx3MpWpaPquJHmnWVH9tg7O0RjVyddYM3CR1Vh4VZPNcMhYwcYZ
FtIV/Ul9o4oUtdOVH3ye4y4GHd/uoDMuzOJw1cVcX8FWaM7YLOlLoXrRttgZ0hwmuFfksJBy43yX
l3yk9szGygUceAPyZyzih6cnbD+V1vbVNzBJXcENha9ra0JMhiEBR8ZKfL4ftt1a2hfX59QGInqD
GMBbtTt7aj0XEmvX8UNHE9M/EH5yLXcOYRypyH1UdenL1gfh8qJdc8GJT7cEIy+pzvlpHAyN2uJ2
418XfkDCDz3bWxCmbkapWzucGp4+A/FhURlDQH3yGIi6WTqehLURsroup6nhaFKv6sJmICTQs+jz
fxdq0zQwMSoJn0pmjrRrvd8v0setoYt8yZH7Qp3NR6MTdyQP0/ZaAXPL4AFT6ZFnkX9GdLdONU0f
5t1MxF2oqYIkAZbQW7uwNGuknFV28tg0gaOrcZUbKYHwvieuH8HPS1x1SjoO5tUkvxJBPdVAP9M3
x9+0+ZUex+Nv8w+bL028r+GimfjOC7TKeqXrLiCFUDIpvCxXQu9VsSFwMCLUztQUoo14/Jy4FS8q
dPZtt2NYRK3IKfrj3ygUIfeMzxAgT/4rSBPfUoWAQXHLjVcUrHGgO3g43GbBjdrfqRmQArJPu8pm
79pl+4txBJkAEgUELtZWurrkzjNZV1YBVobFAoHyfJaRh52L0+3dPFvVyJAqUIyclYKxbNdmVTu0
ktA2wZd0kNVcWFpNeMfbF+k+74r438KWStrB94fYjtVoW/pqPqTqOiEi3i0ZseQH3wOhLE4vw8q6
CANdlBizVZfPrROIaKnXdrBFKt2SW9ch8p3ML1XS2gTy3VTsqcRo0w1wroViEWM/DD9dLFvx+7Dm
wHzqvbpYAVxIS5zekJmTx3+rjlEibY6XNO2KWnuQZtoOiZa+DXMOApZUWklLVYwK1RdBF98coM/7
PLONRwMO73XuSkHgVRK6SmSg4EehCoIYxH6Njfh2mbS5NVDMxkQMXibMlYErj4yDSYwJ14sVPacJ
zKGL0YXsPcf/2xFQNBzrBMNHmjXLxoL7Tddzp6QjYqTT8Z38MgRI29X48JcLLqzW+33wQXmDAay+
FyDQSZs8aDFAmEm3xalGdABXnylv35eCgo9dxxK85budwvKADw5qvDqSK/7Bk1oLVMksHrPB+rxf
jFpzwCkovh0bjbNyfWnGhQPxOLSKmCFy4eAiK3zgQ+Utg1ZO9IcdjYWXclRfr04NkCiJQsMUeaIt
pLRpLzMmVh9yXsyP5Zait8t63IzHV09Eq2YVdvT4E/UVwYX/fUvgqT3/JYyRUCgXKdU7nF0ADZ3U
dno0hXQ5aPPcNobmJ+JnDkGo3UiTYq0h+KbykUAwcq+14CEC4cQiWf7AWRzrd9D/DD2kgSd5zDc9
2Epe/0QhLiteN/edY1IAIYfhZzoUjiLvONdh33DfRg5YyeslBU3V334e/hqofAVCmc73i4Sxpm/1
S4FZw9p4khvtInnb31WSR3kZrVadfux5ETkn0GtQQgWXQawjF/MdRTPeHuZQu1mMRIcgyrqgPhXH
qxqNz1QIfe+4P/9uqi1z4g88ZYdsv73HW8sDXgvcobJvUxHEcoK8V5t/QY80ohjHSA4kxB9S/fvp
l62ihPtEbkl3C3Q8+qzRPrDGVnBLv6iAchv6B9w9V1M7ooVAW2R4uThg9QUR7GroiupL0LPqeDXe
RDIBHM3UOdyuEEAZBKYPd6DJLmAovgQX50TqSFtexPMtnxuvgschbQIZfVKAUo1hRlYpB5r8tdcV
mc+62F/c852021QVDKzaqNSo747CFETx6aXnuxXt17HM7Qjr3HFMh8d7wIe5WsSV3Vmk71Id8KcS
V9ml+9Tv6C3Oq57AM2TmsdWoj6iWhI2Ks5uj66YBowl6UKMnrhyfW3QkiO3rxH5+IvVcCemHKvFP
DAppt8ZnXQU/n+WmtQ11ggck9yRvbAd8Dz56P95jz+efUnopokhLAYz4m5aH7U7s/grrZTCF61lp
2U1sD+YBKJw97kHHDH/txkKAzZWt1zvzkx1H5QxiVLDVlV2NLvJUY0sDmFv0XOReWM2NsJi4ZTsR
D4HikF9B1pmdUJXWqo2K5oZ3FZkyRAgHBhWHb573S8wxyNiEbeqUsAP+YM8aBaF7yAiqB4Z0OYTH
Kj3nWWvu+EQJNrEpse+7sZvh0dAgRanjfXydbK8ugLDsTw5jzouxav9X4blc4ju/pL+c9SFi+LSQ
xF5SgoDrNMLFve51Ye+dB7PO2eUpQ0o8QBXTULtHLtYfZolPh39j3enaOgmNcLDjc0kZUIdj8yxM
HQhkorSDtlNg6CaStZeFlD59xM++k/StHnmALY9+ClmtM4WNLifDoScxt23BsSwJ757Sgdqgog+K
zjLjvQLz83DgumPuF6ATcX/CIqKewpb5HPet8bYSJwAa2LV4mum8dqstwP1jNBKLGPTPWVWnk0oK
WkFpmhiNK88AKAQSHIqWMHBhAzZ/D8YAkZ/+4FGZZ3I33NFs901bqEe38lCHTrc2Z0IsTMi6ulZM
AcGH8s6zjINyO7+UQCjqyKrwPZnFXoWUI+GyvWhsEjiEdyO1SMZPDxaTryHj+0iKNRiZmAJ491tf
QgPAAxzUOGgyPsMwa3D8BDfp2T5+6J1qAWrrOMWaN2csZvv7RdNU11Ci/oOLNMXhmocwp0IQi92n
KnKjUEyLBpgpABkSV62u7LOrY2LJT38CUR28RZZrgsLvt+ihcqwchM2Ghz8Ig0/qN7C3TJbJSdbT
4CuJK9nJMXMJ8uEUWBzoPE3cVZVIsxBEznJwKXTPO+4zDxxOFZrNMAinqcNPebae2+B/I7++rVH/
AusTsxNCR4H44RtNfHTPemRcex2tIKOSfDHXwPQd+NyUwgfPQhyRRg26AlDSYZyAdYkH0taZVyHJ
fYtUqwrfiJRpKTveqj77/9LG7LwXKc8jltvjuUM5vv+Hzvy022sTcgjX5T7CDGGUyW/PW9bxCk6k
26ws6jubEeRKAYzeDMGypLcpgIASUqlGNcySX7qclr/zJkxUM1NOmHJMIAq43kltbbaNP9qxzv5S
aNWAkF8o/2uuVPJ2mj7dKaLgVWKU8+dXkd4v4WxiRHcOtzv1AuFw2iSnaiSasX0s2mmi7Npraszm
qa+a5IaySPazmS6xKj0OO8scYagqAq00knulNhDF5Gzxfpj/liHTQJHLRrNa0HS5eYSoVz7AcQ6l
cymkIwJGNSbnBvf0uuaWgiV3P/Io1C6PpRgTTX2TvgtrKRvfOHGRcaP1LHemVFRpDVlAaxZGI82E
5Ex91EhTuLCF5KjIOup1GC+Rt5z5rnXAVPuap68YT8wGlYZamrwWfIPiBAoK6hQqPow9nMA1EF3G
iuiyOVXjpsk8RgMlrZBHXMs2l1hZgdtC2ci/+QsFmWoUXXtXlYGuEl3tO+jxFoh3WaGFFLjHRv3W
1JlUW05pKFcyf5IojrvJ8OaV+20t1DoPmTa1CTIt2wCFOlHxPP6TLTOuAS3xuYErSGqmU9v0uX9S
Ij9k7W//JWRFjewo6/jFyyjvxZQ0TJTlj72NXcc4i2b3e4UDZVb52HCelJX1G7+/bWxwx/gf6BMf
0bNhMrP/7g89IkttnPRPJE8ATq6Y+A5t3ntPNkUfPu15Fag6sdNTxXeknu6L0jfvCd8R1r8rHDaU
gpB9mH7fzM/nSgL5khax+/n6IGwvS80+/A4vJbnRsSKN7KdzF+ALBjqEhga0kcm8ALNdqBnRwczI
kCQ49N09g1/JENpr1yfBAGF36JL+KDqSfQSY6Wlhhi/CjbAmKVm/aG9cLl6ecByMK5A+4ePePagA
fDLbq62cluId5Uv89bqF8kq1w76whCRZeVsVlDuhs6TCkBwjvp2GjMiZBe6ZlMFyn4EhaUMkhYHF
1EVYjlJPCpmgVutrpb3+OKcf2UTrgdnlyAoXqkCJNllMzCF9ierjRG8S1Y4boleyGB5MOsHvz2xE
qiTkQbfNpLJOcV7U6c8GU+bhDVLyi72ItMJq9cj9Od6lPfTwXqckwAJn0o+266jricj9M+Jn/YNY
0FgHj7ZH/pGJq2WZWjnmRBObN9GuECNa7NrTI+UfQm79aMjCxR9GkAcaIBlh0cOf+f0OEzwBXIfU
buy+iSQz5AoprWkNAt0i7cyMG609DBbiE0Rkx33hLnHZu0l3Pl8DLumZXsaKWqHkMx6a/ErIWfia
9JdNIfk1MvBD0woailv0BB6D6q+txnKSM9rkMeeJYKuPu9UvkvBcnlnMssWXZeey4s/EK003JAjB
2t0xFFXH1H3DxgkA6SuoshXt3+MZcEMByyql0V1OVXfENqmUdAYRf9Fod18T+ktzxt2PIp3JMJZW
0Bz9RD0UqykVJskQ76XQ1auhuuWoxqMAymayVtzg7c0CZ8NZofbNMbYbiAoLgZC5H1pFcIK5IXXA
3MscN7l987G2DnlUFkx+hSOMEiU9I7Paqxd8fPgYCC3D599xurexxzaRAyUOFmdMGDfPLRV2lm+p
19G3jXOBJHOG+A0YmwOJucQdtd3PjHJG0HkizHqkVzEqVcDXtaYO+LR7SMtW5dYwUIlUHZ3Orm9x
rSyAT5pAi4KV5eD/SPTAjBmOq7A9Q+NEkp3OeB44cox90RTaGzT19spM81qOxOuX5UztX3dYj3vp
VxK4dn5U/LfsPJV8IwWTR5y6qWoq5vSRh02txxd3ALjVwd/ij9MUtzG4iKchL8z5hEh3Q5/bV/gf
uX76fD9CWccrKOFkAiARsFBW0tJB3q7IqXmHePgMdY32hd6BwtHtT20rkmc71I5RMvo0yALCux6X
/0KqL4LfZ6BdmJBYO5n0dXQE9A3JBDGK+B4gh8jLOgc8FtZ/MNyvPhRqlHDgGlaGXhz1zmxwH4ji
urf8LTFZfZmwuptiV384pkQqExggxCRG5p6j/frH5AoI2YzPdGW8yawNSAU8q5kYNa6PJtj28sTW
6T6+g1Cz38MLtrdOs8J23KK2UieYLRh5UJLPeYtXJ3pV/5NkWbyG2H6Ve+DAHc75VTRhEGEHRAHn
dNF+NAUt2a/Y3+baA6fzOI7izIF40Rl5LNJgOoA0GgR8SIUxeVmMJZQNmqFFOtGpZLahfIA92HmH
0ZmFdZeyR8MWeFYX4hx9r5jHeTumuoHHoKN1TqCYVJJXqnXKtpUkSh32B9p5tpw9Tbl638BYkXqs
4y7JSTH9So0YcYD7ByON4YY5Hx4zxMLqZZbjrgSAnRX1AjzNF38k9I59QYuQC68o0O63N13Qi6CG
MD38LfN8kyeqqrV9hq9Ru36V7LLtBq7j1zPTwL2rwxUOmN2tqb5Fk/lnCNO78wgRuXiRZjC9oT/y
T2O5yb5PL/chhkdzV+MNPpn6l4oqMR4MK4ynBL5icaFN6P0BJNeXfakjZtrzCGXRk30+L5OY4qQX
t8+qlSKWx1t3FUIp6Y+cy8toK7+Ta/Q9jskBNcOsXN8iZno8a3rfO7G3F95znFV2L53Gn2rK8lkT
r/lfzTeU/RTEjilhaI6nFstdR8PyiiAd0D9ZUwW9HRJRV2VCVx57U4ZdzqDbqNCTHt59IKYyaWTT
+pz5lpVOT/cVIZHU/hLmSZlXRKqJXNinHkXSvGJmHqz22i7xVujlBUNQwv/0E4vB29LeBMUEeRK0
RYhwYvu5EIcrHeDXA86Wlrre4uAofCF2KlmMgjX2CoN2SAOVBmJ2T0yB912fePhdSQ5CiB/U948g
1M+gpKeAP6eLWHMPS12gVlY+82/UGB7CHwntPzT4L3kzNj82jVL6fMqJswBJ+NBLhlPi2GyadfpI
yN8ZYmEHxuM842LFc4EApLEW/ou+rxMs4ijZtzpF88dnEwRFXYDrH9hsUcR023TQGE6tFAuFFdul
TYpJdtRs+QZKpF4L8upGw7DT5Fl9hdG1Db+DbNT+6PVlzSV7dbrRwcx/MWMG7wjLsHYeI7ChC92T
NTNaWMRanxXA6mrHQU7x2yOpNLSomdBPCFuaNjqVFfljBpzIl6Sc/Obr29OJwgREU/N/XtfHXYgA
oWLiQjml61Uhzp0NIfEAZ1gusaEJtSb5+6/WABGSRRMc3pj4+hUZ8WCd+gDSy9hncrCmMr/txUHF
vabhLq8vZp8nWu3J2241pArue0lke3AU930Ef8uIvsN3iXYwadiAEPxU3Ik30QWSQlqE5u4CsI80
FR3EwvkJO5yh6CWOEpUOgnesApR8iIW3tlVP++Nq2oH9F6XyCOTAtxad4+HF07I1dlL6u3xUSbSr
SeXx/3k8BlgxH8HMQKeNya+aMYs+KdHW15ERGjwtKxqJxU2hmGtdy28TIH1MJtt7N7ofqGynCPcz
L3MLadFVsEUo8iObcB4mwubEo6blaa2aQI0RGTBZ/6eFjl633JCGvXbehiTTvui+l5ykzGTXXxBi
E9hVHrq9GDjy39JshAHIalchGVRkwQrlUZpZuEKF0IR4BeTHXfNSQ2EZr62nDKpwz9u65MwoZDjY
9dQv6ApylN94yjRRA0wbg5xLt9kF4EbQOd8an8xy6M6PUvVTfxMq06wg6Q3XPQaxK5fPvJFamL1/
G7iAIDPbetZutoEy9gVBBq8hZ7/RixpZ/8KrN2ZCer3tfTffTcCW/sLWnYKwKubm2crJKYNYgJgp
9zsKnVGqeWVTsar8gutfffI9PxlyC/T4J6bB7sUT8EvZYSQChmmgFh+6/T7srI6FeyBABRz473MO
hdvb2xYjVlkEFYz4ES33RgJ5wtKuHXxLMP+QmrRosGWhpUA9tKxruUJLFs13zCZ2brWNelmj9DAc
1HIVjS/FKaWQ3H+7s8KCltqwb/ytkUNsjouuqTCKpjGTbROFPdb3gcq7p75qFDlAwl7puSINgKYC
KK6fY4sm6JreJLcKE22MidMkiM4Qh/axo3G22c+0Y4xg+U8lj8AKXAu7t/KIdCPgJ+bfQrOUkpVH
WJL8GzCZ1qipmnnLe+OGoDOUCbeR+8M7I1RGxTrxRzK8MoP+wNOoLOHc20E0veG6Rr1iq8zM1jUc
OH4DnXyPpz0ZLNVSROyBJhbpnHNvpKQ52u/yol06f6QDBUbLHMkXGEsZKydL0PTLcJnB+YKo9ZYV
J7ddhkn3h8eLa4NUY2M9nGUw/XxdWuGt+2uX3I/Pr29BW8FQV6Fn6pgtz1QNv2VdYrhum+lOsBzl
FSycl4dizmg1SlThKZvlioUYYIe94YCw4/PdZRU86U6cKKq2Vb55VQgV0f7RsGb957carGyfAuFy
vv36ep6wvaBcuIqPaI0fepuEu49FIsfAibvQJYZiJjpcea4+0IWLc99zFayCOBIChD2R8Ghey4Qd
yorq6ez4mRjxnQpvKDzlYwtmGrWmBpKgZAi4VB1QJwOD45gQinO55o2NZRAzgwcRRU0TcQA1aeMD
b0NIYfhDHkwSw93f+Ldpr7SFjMXfNqS+49eLm52EOi+7DmeukVbTeyNDvDY0mmeLGHUzmBPzSHJw
MBcFCEbU5kQYEA1udqpPFxbDodoFPq/qxFpvNOxgcE7Fu4lWTSOroIXVDERGPLbcA+aWcteHrvtG
455Joi2R3lFBJAemzdY47cgVqtEa0IrASPZUNfTl8NMtZOq61TKZPVi+b2ufF0ESAd0ovA74whSj
Y9f97Ikkkdzzv9bOT1RoSJ41tIlSTxw0iKA2GxrYJ+SHeObeK2clUK68qwCA57aKQ0V9rmjFVhNU
9a46KDvkPVpiTa+4w7JshVLty3KpJ+C4FwhdHgQW4lipMy8aY6n+NMxFfSzamMNgaaOYGYqZ3R54
R9A6Yos4ngjnSOFxCgIk7DGw8iXyARHOkGFLgJZw5dY1F7bItCmEuvWv6iJdKdFWp8dsMZso2R2K
KfyR0URKUd1gkMtMZsUX9nGh7fMlJpCBf5XH+oP14HgStEm5xxMlMn/UChOB8wrRrTMaUIwGy1kS
UPUwE3fvdETTVj4Gv1KSxAXJY1tDz3+HHCEUTWoPKFpQ7XCExIkLwhQ7W0FvvrASGP8PFo20QTqH
D9qrLgsuTizjH1Jdge0DMhVU0dAmynCR/6CdNgS8jFMEUVONRHs6V3H3ZT2be+gZ2Rt0YaY7J8kj
8DbvjBbXkX++4/IjbTxGc/a8jtXJpMaUC9mweh8IJg7TxFEvnM4/qZojPVVc4D0cFsIQRQVBK6B8
fX3fjuQjo4wRNOwHDepaYOiNaZ/D6PMWeXwhNDPTZJJvsTylEs4CCALVh8RoCgv4/+9uRhl6ud8L
a6R0ETGmOX66imfqz6He40EAmXEXF83/kZ5ecph5nX77zAJTVwwItpUJ/p/A3ZIrlCXb2WdrTB+b
h9tFs8g8iOV1mRKaN2OXjnSTCoFpdFli6psJCk+yvl+wfsjU0WUHeORguY7q1SMStZOA+wNoKKio
9naRpdtosvZ1SPJ8UvzBI9dx/DCVy/a/rPDYTwuRe1wZSeZr8k3GgGLhbOkjVNpzpKMAKF55peI9
kyd94g5qwab6qFJoaqECPUEkjEnYwHdWUIPzpxojfZDKX6RMLvLT6XOvhVKjrasrmBgvMbg9BH2P
u/uqEYYGrft5PbGFEfjPU/wokZLK6eO3N8lI3ZdPQftfHLt/XW8YMaMfrQfH12MY0AJVZ4lYmYmH
m32hk7nzV/vn1JZ+GnVth3U5T7jLwKVsd8noejrdK4RmFPXP99cC3yHu9YxzP9g+JQIR59RZLqte
9zky4u3MpItlou1eHfL0NZ/WM5XccdLdBkNNWKWQ24Qc/GUGzd0Cjfi/OrnII2nSlJUzJYe43zQA
oUk6xx5n/kEGcmNUaT0esS3EnJ5SNnDsX8jEMGUDzr2XfLG0S2ZsZgfPSibsOJJvm0GAx/lUrxUT
5+vqIy0gtZbOSSDXROaNgg2cCYJ1JJsMbooE+5IOU/NJCvor5mkRHZslBQyplEJi6llwU9qX3qPA
ZNemIXFVYXSfphTNzEhHKtS0C7w2vTmdBuu4L/hXWEPNFGlutkFA/UeIKTCl4u7QZSGdbMkOVO6Y
r017Vg7cir1Oxwo6CPuUEbGQV7mS9wKym0TgKW5/PQOq38FJ1qKGt98x/lB8V3DcYjp+j455I3EC
Efu25qTkrMnlrVCNUtJ9Rdqi3p96rpVTdiI7sbJjFMWxOIJMuVKPGZGsOohc7CjLLZKOzMCq9IM/
v3bi2BkrJnT3gLrRqmPEIpttMoGVZyhgzoqyNolwh2HcZeTUfU59NEgcTaU91XBIK4YNAf7fFcIC
owQ8puazodwJ/W8MmhMrYKb2rQz1meQLwKrJMgZZdPW6HeO/qfiWhksnH1cPWa+5Vy9T6ohPV8QB
XfHuP0hUseflvkH6JTfprvBU7+DpvSnJjjm54rgbe+AxFGYaKufnrw126QnQwxQxX4Rghg7bMAIH
OXdsbaiB6LmSXdbr5c+RGscrW1+L7bJxTA5XvcTRY2BZBpWwIvGG0tx5UhiTjSecoyaztfrOinfy
welu0BBChmcvjSdKDRJKxm06AOFgdN6QZesYV4GLvqJwBzpsL2nGjvIZASw7f/vrA7hy3pt/lSZ/
pbImlXKgHASpX9VzCu74Hlxx1TMJrgp35P4w6uIg1BpNpltw6qnh8tPW14A1qQ8x4vogVlljhfMG
96CBrB5Ob2HnGohJ1j+3cFfx52+LOzXO+kNVkDd4E3NEobKRUN48k5gFNvmx8fDwQ2os4+mZxP/y
YfNox+lulssIOKqvMQbYqP1bwDhMzly9eZcqh6Fsdyxtq395bXhWqqsyuoYVJN+zQ1POBXFJfDXM
iQA0cfEkOZI28QRwhJfGQrojhZrTMi5zrczCUzKe7N45PlzZYb2lEW7mQkNjoehwX615dIhY+W8A
KK3V2bMhFleWEIIxl6UdPa46NiMwHPJ7lHystZ0gOxkM/EBr9PiaZkurXhE9caxy0VASQePTkVtX
CNwp2rOg6dx1C6WLpsxqg2XWelhnDl64U6AKIg7Ho1NHsJxWegDJPD7j02SMS71Ti/baLZ6ynM5v
i7kUA+Kw117X7t1cCiDnEkQ6oa28sUGqSkUN4SmBCDyZuA9T/P4EJPD92BGw2dhkM+UmLdf+Cz5C
oOKmMOkMhMEZEMutDL0I3jcPMh4GcwCE7gPAQpkx6Moskq1taDMDepsNIjKzYlggZuvubAgOfqk8
KpPP6sSMoobXv6guoZ/tWaomW+KQWXkBlbC9ZzHBlJPKcC5PxQpgumpUcUSWTl5fBvr5QqxL2XXW
XMTffF6CGaciKg3XKhIEnREVkK3ddJiXv3wGzlaTZ2CVlsOcuW7nZK6kXfbvPJYYFBmAjEYHCVOQ
sOzQstEAcewJaOpvTEgy7kU4vZvKoq36q5WknbzD8Q3lryx7vcAUsdDZZfOc3F2olRiiuNkDOSEk
fNnUCnH+zvtb5CZfdBsL/SRq2pjlLVRGDl87shginCO5vn+Pvf4jkFaoPPevTCcQBXVfGNwpVrxX
TAhAQqU1DEnCXnrdX/eJRzMI8Q5r+FK/MnJSYZuofGDNlvkR/nqomAyuLSqbukNJxnXJsz/NMeU7
wollI9vwC6UNP5saQcMaqYS5QwQdM+Gr0qwlFpiCH/5KXvOrd4zCFjGV8F35KhUM+z48EfgOsvMd
6o8HhIGOfOwZUcPxsFPrqt3hIjyU1mWJAw+wIbMPr1xluixicNEI412LJuSDZEu3fiw8MUUR4ClY
ROO2bSF7IRdJrBECyF6xg9VBISWhY1ZizrrkF5+zbGgFrFaWb2fHzTH7EGZjoejqj3wC1DnZweRN
+nWOQkv9L7XlAmGG4QDqJxjoksukFgD69T0odByS7eCC2fHQIcJMYc3pjtgTRM2PQjREIkwPLN6g
Z/Sv61f0Goj18Z32A+SiUHF7fKDNrGQI2NLYBB9TV/RDkBnaaYVWm/5fQQHOdNSn27UcgH/JMfpx
7EmZPPvJvEAJ/8GMBpMObZYMXmfE6d1zJbShxRPPa44QhcorkEEKo/QKrPWeVCVW1bmeRXZEZUOs
8pNYOWvFDp/ifTAmZ9xwpizlOgSxgg+RqhPeeGkSxyHyF1ha1PDc3ird0mCrn2hsvS1xuiCtMx3H
Kfx1vFYGYphY7aN1H3kRxNiAcIsIt7vUgvZ+YphaA8JtN6OsZ/Wn+Fezy1l4MVpTStq7s11k7Jy4
VhoLNqLAR+aKokOwNyUUb4DbLwEXD0o7Xb3HC5vo+zY3ARMAS2jgzzFEYB67ptsFQnIhfCSCQjon
E/J2XawkJmHrbA35Bx2kXSRbw9j9J/FyvW3ukF/Gt5mp6qAFT+qi7QX0F6BjQpdj7QDRg60APoN4
Wm6Xf7ZVZj2pey633h5Qj8+nzUhA+UuENJuUgzWZE/R1t3hsPQgDpGlBFE6iWMMgkboRZpKvFdAJ
8kBtpJd6q5YJ4qog7Z5Az6gqXUNFkngHu+GIrY5cyRnw5UR7YLOd36IeUqgZJMONK/6WloswjNYO
AgA+XMYZ2O75Dr2WN9fnEPABsVENG5DfJikSrP0WF9AHfB2gCK9M3UKnSeoVDwGOYm86NCz6snNa
sw2XMdLutzJlSIZ7iU7seTxIaEGe7m1YdIMaRa5BJBLebnsKbIZgk1xAcQoG7uSYSLttzyx9WDcK
j4fFrTW3c11kuZwiVAnG35DYbmgOj7AM/7PRoNTw4S9EqAwPQ5JMrQ+Ettd2vecuMaJDqeseMkID
ubTDv8+vGap/hlZlxYIT4bJPI7Mxtxo5zver5X0VyBjSt4pdO0xCrM/275ER99PPEt2DEO+Hy7W2
FGG2r/d5xInRXI0an5giG3LlYLDk4N0jdP7kKEETY0rH/9kEFOmhiFotiJQg+lcRlxK5p0Z2OV27
wr/ctFzqTn1F5JaIUJ/vAsPdX6WEiHrHmOGRQMgB7Sr6yKwo3x9I87PFxBQQU2eekOY3YsxJifIt
Hzszg3rWkFjrqEwOC3rf+g+f71Ur71Os8KaSsf8a1Q+RGyIa2fnrAEqGXQr4fMa1ioBal2h2nh5j
BY7H/Iy602KN/r7OVEesCKVvI8m2mHYT+Te5ecQpJsbO9Yqj1a1dK0jlOjpAUV11I8A4KIDlAof9
vCNpeIC6+B0GzXV2YmnY96waMwXoluRZjCAc9bRLeSaR8672WJYS+79HTfWG4+42WxXT+Jxs5isY
zmSW+gBjELUrAVKiZQuZSCg8bKxUXFF7P0/4Pm3RXS3jQvitE0EU0wX3qOm1W0XgCrogMzzV40Tt
9oGGJusXwPyZnkPSvDFtKukOcPkPWZFHYibkZJpJPF9oxWMVCy+nKHcBktyQrKZaO3uqcZvBWvK+
QD8koto2QDNkR2DihBNoSsNJnhVAJiVmkgphYGY/WSOqtMzykAwx2HO4ljmBp4+mLASgfGCCOb+V
ZNeeIh+EdOtYZihcgFnN0Q8E4jVD+GBrxmGA9V3yaRY435qo4PA/uTUi4M/THZwk9Fr97hcRtUsx
BuYXffCeJBO59JQGDa7x0AramMyhtysx+5t9NvJSO6T1E2Nn/SQYY3atKsxidBJZU5LVyQj0S044
vPivyZ2KzJb6haqHYr+jGG3/OQzZQDF/PuQLgbV6aflyjV/6UPCyRzrT8OqGTOcZWDeAKD08spe4
H9GbQLT2WNyOvOVtyxCkQ2gGvvDXsWfEeebCMLSJ0mTZiDlOr/g7+ljrwzzd1bbYO2cV8Tyc2q2d
7uvKy1OUvfXg2t9LrmyfH6/z0JaUULwUI6qNoft5HqX5QKY2bgoNZAhE5UgMA5703RGPtZSLN+Sv
JAp1VYhhTMZv9rnrd4QSRkPX34nF4eghshU5ECm9G+fc3w9/Vx1vx9bu3pY2AtZ5PWfTOVHiqOa8
Wo6norWodvAZZXOcILKbWrcX2kTUzFmuPGp9kpLT+w3Vu2CehBpIeVtiHN+K2yZbyWq1e9bykJQo
MuAXzYnUYXlsfrCuRdsARBz2pGVBPHY9roXCDWdQkW3AyV/gKXDK2fdIv5wxMLH70jsnLwTlWoTv
gWCjtaXWRwvHTBxlTwRJloVjPIHnc+5c44U7B6se6PkYG17RoMRb0WFWL5HVh4D1f+NVs1V8FrNK
SOf9kdcD40VNcfvWlU+6/jGrdM9+jFn7NztkJtOcuOyc0Aa9eKiwpkkd/MSZGwNE5Hxvu/Mmas+E
3cf7odT0ZhG6Io50h7C2fEwrkEYpPAF/drwkHPUth0zY7x/iGNG6Q2j0yqinMe/1tXVj1HvdSaMD
Uf9Nl340FSFVUmG8KKaKefjd4OswmxzU3sZd9eEds2ISCnKQQka4H027I8NGh6jYZiYzKFy2q/vJ
XWv3GgalaBNWx5a9yV84o6LZd/Q4WzQNQVxgQhr0392VXiW2DGxWePpXleoEpRHdmLxmTveF/Cd0
G3lj5FoSIu5WQ1iEJ29KLdtI2J73ou29QcSqdxHiaIxDfqoCicMrYy3FpX1191rkS9qVkW8YbG6E
iVwN9mgWmfRWkL3uWqIP1sSNDwTJx2x5GQhoGmSNWjqGPIg22NEsTcEox2+UotArO3uB715TTsVR
uLS9UdqE1NWDAc3ecFy0RsdZw5K+AUrG5Jqq7VWETkSoIT3SkL79QUWI1YB7SCDVYTOMFKKpTAld
tGH63JgXMoWBiGXQYncArgTOZ8B5Zmsvm1uyNfypMSvJuZZ5YnEl5u/Jybbp0Id8LZWd0pDaRghv
c8sGhG1oIe5gTV4ejk5n9f9yFRGh1nl9ksQa18lbur40PVOEjwba626xoRF7SqMQkXorWUvriUPs
E3wGAVv4QHwbWJUZbuvPa9638E9PpOnikcOzKvXZBcScDouhHl/aklT+abs/Vcfrb3QRADw+vRF/
Bzff9t1XWa6ECFbPNVkdYho0tGoQfZw7TiUugYYbP1HpBhHvaAIBp3EvdgquU3B+sqBwjhCPfcgn
ObTuYg265SW0vCjC+wZ4ZbjxAjA0FG53sKGh/f002+T5R5are7bw+qUqXqCZ9iOJmHfBQLIO8U5k
jTeAEMf4oHOHZm9wiQ+mmQVT3/EtYPY2DRsOfYiWogRyxkq4/L/jrXgjbwLItw/CwRXPFHSV/O/y
7X6jc5oMt9Z+ynXv7eP6EHKRH5T61F95yygq/iBmpmqrQQ6L6aSmNyeqYkM4F1o4OBdQIfMlKHqj
RW3FChsBR32uCvQUSCoZNf6UzGRAri945fjtPR7iXEBvywBR8xXNQU1UaBW3tFtvMgSaovdK22D9
xNlwyix5AAiqkLOkJZan08qzbrLU0eJFQB+jzoymjx2/4oKJ+IRvO8SHgKm/FvOiBaXoarHti3JZ
XRBBPhUnPCIALldLKwRxbG11+2IxRX8pMfnMAD+3FOOY17PdPXuLWoYQpIDkZFZfyRcFea2D5CzA
2v+XG69TdprRX4Re8XMRgMrgKhHSEh38cAhs+X+lOtsd0vsVqfp0H4l5Bcp0Z+Q40NZvoLuEeKWV
7bry5l2DQm93IgqUXtBBccbKc6vSLFFVi15hST7r/nImIELXKeRrGUZXR3QI6KTk/jFEuojd0sfb
H27cuf2xuKvsVsWufRw1likAQnwPwXLJJFKJqUwz4PXVnS2Xg22+OZP7zlo+6D+RYMu3+EindPil
cJSOGp2WaLf+dEmfdiazx8nC+O7T5H1e2TudvBiu3RHqlMG0YiDE9GxWdLD0UXGyYMnBV0IKuLBM
1IFFRtw/Dh9ayYyTE3gAPa1ZUnm9kcMp9m/xdyHUhR+9YjN2Vm4+8jmvF8vNotrPraIZKYS5tZ/n
VwL39GfLnJiTKQqxMOLeSe6BFWePUyMJDBejYwQ0K9jMvIwnEEJUjMJGU3xAcV5LPQIh6iyMsk6z
P0nL3Z7hvUKPPKyTgnEKXilEPX335Jt1h0b5leqe0KGlwFVXr5+Bg43to0mLx5dyxdN9bJnE9OM3
4ZoKjYbz3VUGECNIhyHPzJChlc4itO1c49yPIjsjZw+ERxGcHcGoU76C3fyRcp7g0f1lRk2svpqP
eLiTC1AsUQaVr3jTFr7mBCVAGM8trvXR/fwiWKRP6UJ/qt8Hz9B5bRJHJJWJgaedK8uU9rxP0XQ6
1a3tdXkZzh+yzfj2bD8lwYCvWHMe34zyUlQ3ZcYitjEQPC9UbHi3biVrpnViA0dxheRsymVgZn/J
gRxy22zzrXpQp92x//SCY6RDwZ7fmD3aV/+vmoT1IrAiEfXNFNuYbQ//SzGa6FG6kQFMyOJqES73
GAEOnJlLRkgwEvSxWHJ6D+rgcpRjyu4nCmidXtwJ5BcURQkl/v0pcEfJ7lVTxtKCbIw155+qPuT5
NS4kbmb0h6ydoRFPByovU3vJTrKObgOoiNjb7maDi5+8Lu9S61nBZtVmmpr9ThhLTsIOWtbArQKA
lx1HvP0aOlPU/iQjioaylZxP6P+4U/RLriwitOOmfMYo9hWph6tkvJZweyqhMITrO8bMJSJeS2q3
127zSjsdO3b9l/CKyIOjZdof512zQZE7HbPUeiOLxRH3XN5elhoPxhqvYuG7GKIJB9+9id9xwgYs
EZL4i9mxop8REJOKnCTtekXruvhgzuS0bKKSE1XrKZEiOM59TodY8N1vS/baf/PsL8XjgvCSbTGF
oXTTjMnkUcE2GA4QK5FVPh16wF1b0O+a/zM1dyXktT720+7SfLdyKXUupVvI6rkwvJiXn/ezlkYp
piXpGC71w09KsaSN+kFv8IRWTXAhROb/7Mjav8SZtY6AIzW2/wKt2EkMqRw1F+CNCpFn+cR0Y5c9
Kelg0YRZiKrdA38XH+BeOh5jmMyep4yK7o4b20bkzjdHwgBdjGKVAwEqIqApK+4J4tlx8DcHbmSk
7YArCUtN4WSEBJkmDODkifaJXcI/OXyoYOOswLgCT9eetyNfrSsh2NfaB55ifnecZSopH2nUzhtb
DNgvd9Mpo0lJgX/aSQ/XaRaQKkcEyDjC8DOr7e9RHnyQeiz0Bss9PUQzMMLu0txiIQq7hVCI/81r
FcywcwU+9z30nAOuH4FF4EmzVrOy4/mlMNJluVBsn2eynuh4nrImIrPI44xrCnDpjS39yoyno6BP
6e3iM1Zrtv5m+UXPYD5QwGwIShJpoyYoKzCvCHOw9SeeusMlweOuVlmGimNfpR7iZeUXF7zk7emf
zu8mBfDsMfrXZjG4DD3RWUZW8tMmTye7SIiFJCdBP1EBGKkYvI1qJW4hq+Uj1OOu5AmnVEFMPV6x
xvU1eksM/WC7V7i665Ev2L5U025ppKngsPgWS85Sgf4I34ddWLURxawxd4zjIRodZb9IJWdip6Qq
ay7Her0QQVPBcxkKftGKN+FT8B/GEQVFL0G0Vt7UPgnLxAoIpoFfqZCBuejuHjm/eo9fRPvXAoA7
VYXJcAv3onBSTlV5O0uhiKc5ZBV7eqmKE29PzYESNA4iANNL0hbKbWphstRify19WHsk/Q4Ojty2
DyyPy/uGI2L7PJAa7GaXZFz/FjFXMwmGQbypUMtyv5jEisC+ypiUamG4oFnS2Zcc0EcquQcSqX+e
/RBDdJC3IRdiE/soCiyGBBn66gV3o43Y7BgX23pFhFAZx/1XmhHL0H3/pwmeqtqXNLbPvdnJ1Y9V
iRLiGeIWKWzvWSSBhPbPmbpBOAdxD6I7YlCpSqtAHmlaABRqQSaK9b+LCOCC3Xdk8jYaEbPkzIqy
CnOv2mdkhg1SGbcNf9+tXDw8MPVSlHFY5eQ4eOzuhQsxG/CGlZcqFTZ3DsJ2NHOM23iPV6Jxsj3r
xst+EEC92usr0XBsclBooGB1kf89UhiU0MZGUnDQIghYF4BUw5sWh9yURY/DOaWU4EfKrL3y0t3e
Tj6+bv6cuwQTbqrby02Md072OstMH7dAxSVNMiGd1IciqtIZ5Pp9sq2xc1trTYOGE7OPnDCs+VfO
7mkN9ntUDuLcetig38JKodSEe9ujkjo69YAwYdTyLowGv4nsO4FJi7Q4HI39/GmZljMwPK85W1Cn
58brnKUf7bAQKgKSIZaykzH6K2Ug9nN+GdTvk92hTlXzrsF7tSQxn/DjhUVh3wNxh+qDMG1USM2P
6d3pvobXvU0URf9LRxRbq+iFK+MTrHe50qw6HYf1hNMNR8gmnM6QWoJioigu7j55gsqdotl8eVgX
kXaXLCPECAZf3ztsyCNTSBra30x/px30mNAKwkFs2+gcYEo5L53WLsqDJNA36vtbH/LvF3fh6V+I
LYOP8eVx8ZcIifiJ/mQjZhHdXCxBYVhp5eCGK+1RsNklBS7R8v3F46puWYdHBIIcDIMwmz+MYis0
KIIBHncWHouEnKWiRbOhoktHfuOT22azsi4RZSYi0K73QTBLLsjbmCMSs/q1SLkgWTuJKHOsGK5A
X/UJD6mXvorHdd6208zaVLCOqpv3HnaHFKncWvbaCbOCVKkC1f9tAGYntWWaPzT6TEjLUEA3Q6u5
uNePl2zcJGexnLhDUHN18GtFvjMMzp/6hFFlkuiI0pgllaOw28kRzNLk/rgOOKNwIdxcJSc4hgGF
ja2zKnu7+2aWAb8XNgjSHdaas68NGXUZ/UTR3eyhS0rNVKvEfKCwLwN9LfFJ4EfmJqxNh4GgqMzV
TD7bIgeSIqclmUPQocFWsGadg2i1th/BPjrPcHvjf49gBCQB5ql7Rb8uyUeelEk1yo3rTXoHJw3F
CIkaJRbYFyZJGNczPMDz+rIM3FtWe7bG8QGmdT4ZQ1Trxis/VpTzGpoot6rZdkHNeEzQYIFFwM0s
VApqil67gAfrfA/I4K7B3UqIX8rmgRCgkdY0HBYhP56yLMfJ81Od8T/HcMbaHgI+TV2Y1EArDy7Z
SMNOnWURE0heU41cXeV0MwLcc4QLvhGvjq8T10xAkond/wN2doyd1oVwxJGMuyB7+1iRGDABHlYQ
ZEA8umDWBZ7CBy2EAhzJTVykj5ZrjedV6ULioHsWO5XxUgix1+EgtH1un7rWOYjnQqi5ki9A2zE3
3Kpj0c+QBIM3ntN0jZzmu1AgjN1sfFM/rYTZvLdsc0P2hkj+YT8Zs5bndeiKBA+UC+486oypb72v
zRXzkxLAWMDp+174PAWbunKHvAAuwYIDwwlbsyrkIAKdIdGWv2rULmjk3AAAoEuo49Bh44MrVmxf
jbUBqrkqTdLcr0lXypM9iESVOlpxPiYxQHvE4Q658wNZkWF7M1DL+glaIYhfM2BWvepTqwNWrUhM
DooEqrLSQrjJglP6UHRz5yTuw3w/az8qdWSOjld0TzszB6XJM2ppyfL2oIuzbnT0C6BjVrzJH55G
qjz+k3EmE6jKAf9OuOziXSryuNGmoLzvcNDoq5OZGwOjpp1jGycosu2F/s7pjvznbvCtRGyZ+jto
xFDv0rPL7JKtBKW5v9b+xFnmvzW8v7rLTDIHQmJe+G5NlSiRxS2EyPoI670/hfkhrPZzP7Y9XLwC
HlRzjh5PXmJonIXYG6f7bsoK+Xwn3X7Y9Gy1cngVNS/LKbL24Wf+grpaCb8QfBFQxbWFQlZnRW8j
qUdar9R5pzfi9m6pPXNhnf6z/Ka2kmCI6fw0bGa43zhnpFG16kGKYpNZIvxY+KgV6okLQ79GRMD3
3Wj7RKpl7qWhzMYBl861Cymq8n+ZXqVsIGWuOJE0pdZpXsO34tpCZnUGffcZVtXIErrKxK/Xt9cF
McAaNYLr1Nzxbz1VShpbLMHM/Mn/V1bxjVQrWDoXV4iWpOrMZ8PbaC771mxD4+XSLsAxYDlQjjJ9
Pjm15UVNMRYjNdJiZijdCvldYWo1GdJ7NCHzmgqjN8rg5ELX1oyRFKDxfYghhzjXSMplXVL/NV3p
txjM2Ks0oKjE+jQhhSeK7ffCgDWR68+thKed/2ckmHgvWYfepXg1ZSpN+3ft6i5dlS9ifuC+1gg6
IoPFak+1sLX4KjCbJjB7pJvOZsuzi44sM5zr5+l7uJ9BHW9xyNDrAUm+CdGJRi5nhHbQDBzO/NDS
h9g9P493tJ4KQERpB8vjoxMwLgP3SINeGlij9nwJbQfWQfat0KIYVHR2kH/7u0h20BegvXHqhAJC
lOIVIOx8PDyHwgYBNydm2/lNRIad8+6JN9tq4kkpMdFKBirPeQKJleWkzuFrtmGmiW84czRRzYDK
mPFvrpEwBBXP6JlnLKAL02rKLNTjI50bi7hKpgwu+g+dlz2v8C1jJDHoSEDhNEe4OahT4ZuFxk3r
Jli2du4jD5zW37oGz99mdeGsHwIPb/xQY4gNYHANhqUGMSeZ86OKim9/adavhLBrWwjY/b/m7zfO
jajAbPBi29oU+zcP5xgGkUeGQk9UeeR+hPOoX3uZqUi78bR17y+chaCowPFLmSXPgbsn9INv3zp7
SYlSXUi6ObBU2aCUnfR31U/Tck1cssz6aG/MCr7txafLmOSkVYTn+/RU/g817VZm1z9uCjfUh+PL
AjR9dMr+sQvDaEmA0N0Zy6oPlYT3OxSlIk5a2TVbSEzk5sAbjyN9YBxdHgLSDQtMjRL1hdgSx4Y6
Q92bSyGPFzHIWputCS5gveTwWoE8/7u1L5PwEW//zpEFiu3VySthVPM0gtCKYvq81mZxcFckHKWx
ZYK+bZHz3E89SKhyuG3CyKDfvjnUVGkrPy/D6flRyW7lWElIPJyItgnh9osw1YWR4Z1hMf0DkZpX
5L/5Cku5bsyf8a4bNQRlPIkfpqfXSMOqDP5d+oJzB4PH7zAuN+n7vKDjbrAdQgcJtPb3Byp5iZEV
a9YxPvXqgQgak9gfXrXFjjgH/YJoMV3HhzF8jU/pv11r9LDLjTwJpSLbmgKdwwF2HS1Fl3NLjR7Z
4PZ5l1iCvw7ra+/0Hdi2QVi+tlZRTt8drzronitd0cf6Smy0wVWCY1wqaumzYVIGL89/kREc+VKS
4v3aaFXBZFlIYcmFBxh3168eDM2y667dEqYamBfseD2G9DgsBMb65w/K+3ug/VH+pRX2DI4E5LE2
V1WfhernS7ih7lcFxDmIw/7fUwwkXVFfI/jKhyyOIqLhwIESGmwTjATd4Ojy3psCkg9uDH4UmbzF
kcZhWYyLMMrm7/eaG4IgqDqSjXQ4B8oCv4VMfkYqBHJMxgAXUGLlDl4mfOBX4gpraAVcHbjae21c
tedERjt+Eu4t/IW8keUpvGMGnP9BWJiqEsvWG0DW8vCvpvbIjp1pBpQh4fhv4P4yyrVihG7MaKbR
auV45MO/dy6SQsM62E9gOEwvOkxxVan/ptLSuuuaZ8VtF0YcOWEDLrDAU0E0emJKmT1o8uH9HfmL
2FmxbRYfBqYGy/BqpXotMge7V45/AA3BwbblyFOBv6E+Z3jXeCDV4NslhMQPB29vDWvxluCl29tc
wO83uqGxHHPJR+m+dBXErPqe/pie4Bl6aVeDYCwN5i12rc+xdQERDeAVUJ5/LQEtyTV1TJQNUIG1
KOO3BGQJokMxBDU3RJ5h3lYuGnLnAT6KUAlgmX3pQvfFhRGf2qxNpQo6BWwMBIw+YrF1Qs3s8kRF
9QHZ2da0zGZVfTL9mV0NvYZjmxUpxv6/HvwyP2Aa2VXDzYdTQXvVtW6ll1ckjljJtqeEpG+zOSBL
rzwpbvtChrDkNgpx3jgx2q4bTXBQgmJMGNAhkqUxMI3fIH8gDUsLHjdXcdm0vUGybYkTBFUQWkGV
EgbuUpNaLRMCaOOGQSCW8SlZkWXK8kQu9uDR5FWvmIWR6duL0BSEX/ymmXZ8ntPBEi7VHTe2Q7lk
FKCByEIY6B26wc0DrPPCILUifrxqmFWI6b4Gr2YINcVt0KIfZgdzvNOya0d4Axf54xNkDWwAQKBB
easrnxYYrIPDzlRgmd96mqjxqPi/pQA7rHmm9mtBhMii2gFascbDhgXvIaZ+JkCxSghvkgd+iy/s
18GjvCMitXOfLFV1mcfxB/8UwzOTnOVdabM8uLsYdUNaMvrQS/iUNgUkonw9LxVZckbtrCAt4HZn
jm47sTPteiIWjheZrVN8dDNDTIrXwNq6jb/NAA9Ss7EL8gbgNQ19i+PPwzW2YIsgTOozffbCjniz
LFfIrAnYIpOZRRLgb8Nn/OTu6+0dJOf4H+6ssBr/6yYVb8WWFxsbp0BTK7Q6YeUAWYeV1OSafQJv
W/rZ0hKU+fT/MHWCZF4Q0xpUBtDEFMI/v4Bc23nfIq0+EJpD9r86X83QT/fhEuHApiTWwIzqXlyx
92BGzywyWTxpM4xr9S6XupCkO17xKIlol+j17p/4bVUeMGwimyy2YtyvbxGhdfKAApL4FbMdUL/c
RwEUO25hRnbQKPDm5vUBKJWTn1eqeCVcMbT0FNJLnxZJ/lulxS8ognVDZ+/Cv9W4iWwnUM5WD9R8
3zthAoklRAmvAEmm8js0ayfC8jGUPXueDT6nUg5ekWdlOp3IjPk8z+XV747nRpnR2g1/qBDp6VqW
YHEjbZXMF4ehOI4b9Qr87wy2HQALA45HVmBDdKVeKibg9uBmMDi83RsRDls6xATWQ0/71jNgH2g/
z0gHtB60c5vF4e+6U7SC2Jv08iFOBdLp39mx05f4iOLaS/yf0OP6uw7gP58h7Tbx38MdJAE+stWq
FKjCl683l6lrc2mN31oEP29RFH9bEt+IcLTacicfVUKPHUCsUtLfWxTntKFSx08o+9FxF8xKhWbc
eP0I9p4PeD+m8XxhJENbxzhUjPS0a6DMS1P9e6BRwdBYDnZfvxHJZ2rSxcLfeCz3T+hyXdpJeun2
Ev/wzX0MfJjHFMuaWJw87NmLACuZsDDkpjAOh+64GQEreQh8bNiSkT9jhxMFxKADwagVEpQSJIzz
+PO+Lj60/z1CmX15oMNZVx97HO2CIMaDy0SqPpok5lvcKp+P6Q13TU+cUKL19FCTWj4hA995H5FS
lVzKyLv/ltduXcVITcT+ywdGGXL4Bd/nivwkNAuHumfXRbfsyq3inOJ7+psQKt7kShJe72KXZ3LT
4Llg4786p4P+f9AOXWpFn+C2T1ExK7+c8duj7yq+TXeGyjaGuNDx3u6Ej+cRx0SminZIXeo9SMED
eyArOE140mgb/UZuXjjrq9liTBJXXbBVCE0mJyxyrjzF5DjphpzVgPz10B3WsA762kI4Rd/ad6tN
FAfcjpecig+J34yxQtcD4J/brNJtokmlYMiuwcbUjoZBGp30uCenE3A/jJE9N1Gt0dkV0104qvlF
l35+JFb4f4EkW5UtZNTKQm5wVJVSKqACRf/hhV/OgKUmoYmbrhCRhEcouw0E/Fo6bi63e0ikUc4T
QinMdpMJudqHn3eEbkSSJ6tum4C3a34j1iLI1tG99dvj5Rn/rWUs1ZxeNMGZZMHua57/PvbEmXLi
OMsjM//GBFFIWD5r5Bpw0l8xA3Q/QXmXjHwtOpHoxvBJ5F4wxxhyObnB9DX/uCeoKOwSZz2VOS7h
zUIN1EKgkEMSpuroKFD27yJExfXG8MqWTV72KJ2zt+v0hGJYWfNoog5qtnUr0fdYDgOf91cJQYWa
suaWdtD7ln1oSzK3LTHo9G2F06cFWIC2P1gk1BRSVSgIK9RZ5TiNXCNc4jKEKDCt0eUvxqi/qxP+
ixHkaC99gZNKRERkCH48jLNWOwhICJWmnw8MWgO67f1XqG6Nw0TL2Hr1kHKhsExBT8DqYQeZ5JNE
0MBayqkbkIhKXiB+n614bq90M19zKPyizthEltDgFRfKaeekS+yUlDqZejn01d87hAIl7cFrlkY3
uOPcN8wTPMdYoSoD4ov0WVFYNgE2B1K3UAbYMYFe6L7V1F4hUASFTjkPpJU9kdjcfZbApTbWfbyr
TcF4JYyis4BDmMLjD1c9mhcdSEtNQGhdwQ56zBtW3vjpB9EdzjKoGm3i4kInYW/Z9dTHUAn2e0Eb
D5O28ZVWH3tn/ycBqF+DALCNWkQRnBo3pB1BqgY/BFUEQ+uPMw3aURe7dfSBLqboNCOs1P6NHcSi
Fh1LNngZIxO3ApDb+KR7BgF2YmeKXKXWtphT6tFdWTN0Hel+2R3EyCHcmSqIy3qoURSONQUYAVrd
xd1CNGZCNUJP4QpLk4ohqdgPZYBcxdzshv/XmkjOUdodckMLLNwdW+pn/bEKet/6CtDYANvz/Yb+
GoJnMwycBWnyhmcB/8A5Hfu6y5KIlHRKautX5WbUcW17MsqKgElacttNhWA7WYikBKOLRlNx1HEu
7Xm2r4rKpbQO9w889nfVN06bPq548hhYkTFCK8P8WHmG3mkTNJ6fvkfaGfcfm15E/v4EIte82t28
zXvUKV09nJh6G83OxwAaG8GuIthFj4bIZuFQ3O7aMGSOKnASU4aGcnZ4aCWD12c1LCIrcsz2Hx8l
swgKrJYJ7TRHdVQXFS3+tZUyCF/V2ze9o1a5eN2KRPfMdk7WIexi3D16lMtRThAmbJLV9GFTj7PT
GRcaixkrvwTaWR0dpGwI2D4x4gIwS2WYknC2J5JoNJwG4WZmH2DFxZAv+rBpPkwTlPmGM5eclLdO
CU2dAUzvtwBK9C1OFYicQ7P2JCc5flcPCIhs2qHS5mJ0lBc2tQm/JqWYqvGytXBmlidsMzeBRFd9
w6wzLH+2mC6bhRrFc76qBi13+C08sxzkHImFUG/SyG8SYT3DOBI3sTQ9q36kL8hl0UhRFUCzPW+7
B3R8YeN/QgAzyZAyqGssxLlocphMv5VYk5ViLf4hStYnUiEnNusk2g6tGPkJhNWh69Qqe3N6IcxU
cIrIOa0pzDKxjOB5e6Nttfp1WldP+FGay2IOpSqlV/zhGe4muqHSEcfxGTMtBWlp9eeJWbWS/w1U
x0fRXPHhrJm8Ch/YJxKcDsHbqL06tIXLl99T8HXD89sLQ4At5BnB3KldltZU1YsVr9QIaniIRMmw
rkj/J/y03faR0L0nimUY63H/2IO5vjgvlEopKql6W79QiS/YxlStNESyOFS2Mo4x5s9qERwuwsEW
xVIvvTKy5eX8tSUHy1u04crv00z8YtdUJ/B8wn9zDL/bCn1kCuV6qOncxfQ8cVYEQ1MN7yfX9kVq
OjfVJVmJkJXIqH+uUpibh6EPOqhusfxMTLSHD0zwERI38tcu4cFIvvHR43/HgS3ZYnYf/HBl2Dau
bVgE3CrVVSO6JSe4Yetmn9SfzFwbz5TTYj0zDf5CCGvSyl0nisjKNm/wNLjvpYG0BWWiYjT1h2G9
KCBFza46cD9O+kgx40oL5swqF4rDO69HNFDzMxdelunj7UvMTUg+N/15Uf3FWL5DytfWZb0l7PNh
mVtqRlnQpOn1qBb/nQzTYYqpfn1B+CKdysek/9hOzwpPdt/cmuWEbuRYty9yeV+mLIqWFuJ9GaA2
CjRn5GCIK50TgmJpyCr+t0jlY7sBB8CscQ+gsydCjzOPI+gyY85aHpbUJT/M9cuoVz9Am5/fciSP
dd32ng9IzOlLavBLWnnFx25LL4Y+eyBdzTWJClfY3KeTOow/O96VDHM3zdfIn0hG71orsAchIJ8V
PKyKOSSEeT0REhZGW0JTaLuM7eU0abAtESifwgvR8II2HNqkJn/7JV8OfdzDtN9ryyo/cyeB7xta
iXD+uj2RDlAagNRjYL99hcBcDENJ2f5WnEupK9tKCGWsVjFOcal+GpGe0YTYikXqQuN31K6KnfpT
NfK6pcVXyPnCIiQKX/L0P3Cr0kW6U1ac1C+Ykk8xbMKC55aTwvXQgefChaYzq0xrorSdepyT6/50
NcwvTqV33wgZPm2e0Utj3zKLNMGs6cNMrqxUFne69T8y18oyOKQVnIUZwi8RjqonVTMbNTWZRhvW
oo0bR8X+abis3/KTUTEeKJuFtBwt249yeiycztBbuEUy9ME7/KfrGGEaaSTVKDUUH7UcSZo8HjT6
IDpQ7NeIfF9m/ABvc2DQ5zLP4+0BBI8IxxJMSu5fVPITNq8cuTiDp5MKyykde2SIgLWUvHzPTuXn
zbtScIoTp2QKdIVerB3apu5H+xPIABWxl+pxc3L5r1isecTuFtdmLeSriaBAp/5ecPmr19ntgCSK
/bNaKd7rGTM4KOTgNyYZm9z5vPiimyLqFRMhsWoJVNX+SfVIG1SMVhrG3k0wMw5uQnlD1B33CptE
+/NM6qqTOKgVrOCz/Lh8ETjaZ0SPjpF9G1V92IHVOGwhCldgMtx7WtKUAo9J1BaFB1/WJKTFgxIg
p4TvOElSWFxNT7WyIYKB3bo2GOy7HGRijVDOfSzx6ZpLVoc1EThwIphqb4Giik08FwGDDKaKfJ9i
26ocekpys8wXaJMz3lXEJ5llChZXmXzpBRr83/QMqIvn32daGOgXFM/18urIYtHDsm5dI9h+Nhqu
HaXSyT7DivjcTQFbSdWh9/El1d8Voec+DlAFxKBN6DqKeZx3Ab9yY1UXJYD3kWuxdfA6dAdQ/N9C
P2PWkMQvnXgoO1zm6UBvmGPzvfVPNH/03QvOwQDmV8Et9ZTQWgkb7Fu/yy194T397hUphq6Y/XKE
LtGP+2XBj4oh0geZQxoAX6e6h6eFyLiLodnmHQw0UAsfcuh47/adJ1P5CYhAlHteteBRj+iCswNO
DgIkg7jaKjLP2ohqQlEZneWERafLKmo5lm/OXCqoSpWD5U+rvCXWnzFCNv9Oyb/TBUkaW4Z7WcfC
uDeBf5mGlsADxekUyFSlFFJ7ZMuI8tKDZxg8DlW9WUXyl0WWjSbt+LwFwLOe2xhtbfpOlHcdjpMv
0m2/KTqQhHTwhwuZiDgyG/n/hCnJUR05OhyxDrEMhKxCzY9MqXjaYKxIwQgJIQTox8Qy/n7jKvHA
YMeOnmlS3oEiq6yF+uPlQ5dkqcwpJWhGew2/s7Pq4KFOfpxeo8bKw8c8h0hCwDdJkfdmD8ub4Xh2
zbkZu/1Qhgf/XtwjjU3UbN6elg7C8BWiATrGGkN3zReF/ThpAGwWsB7D9VD4dCwmA53HH5cGYAta
MHMfI0EimzohH5+9Ka/OAYGXBn8NFLjmErR6gcR5cRmXLnnXlvuPXHPTR1SWdZFIe4sHodDVgug9
LdNqmstAwd44MePoJrGtlfFV2kKlEJ8QFEyAO5jNb5iUL0FY9EJtIdHyhBeR3YJVBvtAile8ImLo
gbh7o/MuFtAhfXeueC3HdRr/L4N3FkJHr7Ex3y0YNsvAMK7CLTFT6BABrbV7oVfVVqPourcY7Nfh
bhSHEvp7hd+e8bIfMaL37x/cla8wfaAQMPE784+tIBXdK71DLcPGF934mMdgxp0XQD3LTiVMLsED
ZtizBKO3H+Xy6FbBWm4okV1i2yHVxw4BD1P0l0g1Wl+Fpzv1wGArFvm7KHKABqLN5uKc66qcCBXb
noDO/XBWU8nAxH+7JiYZUfqlmLU9yS3YwRQ/9tofM5HRvEypTe4rI69Fs90J0ahujxUK1p9n+KwK
7OvkU7MBe34aJBNc+Lwrw1VNERp7JTCsrh83T3frE405P6/8ZHMliuirBT+AnF8VqhYkxG6t0ym0
MpeFKsDs3evggrzY5CPJziX3SrOu8cIf7kpHZasn8jULQnYUnA7UOlrXsn3gwoinJabhTQssAU4G
qubFzVmrsWsYVNqj3OHi93RXqZ/gKBcp+hsxlyqB9C/ucLObuaiT8SvO6lYXJIyfPcke7zwe2Yey
MdMVppRvMDl/SNFt2ZfiiXRAcFK2IymFmiZ7ONpokg1qJP8WPYErDa4MyJK03xdmk89GOUZwFK1J
1+TaciFkA19paRFoapl45U1GQvlFTkzWNxnXgegtZ9ci3u0dipb8+iZT9NLGxtBRmqoNUyNfxtaa
7F1sccHkJ566yvF/f7OMmbEUy0gPTkg7W/Vf0Uy3eXF5sHQN9xmayQEjMKvikh3lWY2w8MnB/Sql
42ixE+YkTMp1SH5vf9WG2MlUk+xyi/La4creRwFLn62p63tyxt3rLYOKJY7yaHxwCg7FtCI4L10e
+33Uv4pe0oJeBSEHbBUenFlv9YxvEXHEmxSe5x9GWFXEiWebvT+3Gx/jy3gZYaq335uph+Vy6H8l
voIipiz24BcSY8XOSgtI+KzLtWIDBn23ijYOh4V0zs3XAQLcDk6QayF7KZWJ2XYuNIzq6/4qPkqB
Wi9umY6+rzZF9/zRytAE0n7+jiKOpxyLD11bPPvEDgPZrt5QizybbI5uCCpu3rRZHuqKfElKXvWw
wL+1eudQXfMFhnFArmeX7i/8th/DvTQAB4Ngysp+7QMHorEvZqQs9S3cKD2hTTmIvMLvjVL8m8ym
h72fjkAZggOCmPIpb3CmMK8IhOs+M7B9RGkAYiI3xrCTWMRUVd7Daj+OQs11SY4wzrl4oOPYgN66
51KMzIwOjVKY1nye9FDmydptFljHMiZrHbS/P6IlBPQ91k//kLoIND6u+gCdBE1Z9Pf1opVyiPbj
HqeEHaK7NDQ4tUhT4pXHAMfhpbltCAEjz6AIBP4DPMxIy5aPUXW1SWoodi3pwCtOhR/y9Gi7UnsX
4qnh7DrpmuD7H5QmIsJln8GLBMfhH/pdgNLxpqAwRW48hx4uQxmS69uWMAZlrBKDhDce+Z64AWg2
E1wEQisaaX5WE0u0NnfDoBo6rPq87P9DmX3te6Yg1tuZvyJe7aHA/0b4JDPi7tyjA12vaKCXRGVR
E5FxjEjx5fWgB2nzic8qtjGB3pWBGulqki5EUjFf28/Dfb9DJgDi8wN3OIZ8AQZlucgmqXlUPiGc
4DSJvXVQz+SPGBD94UCedOP1z4TDWtF9+VdObEHNhaBUSphAuIXFi0J/CNxWMBg+Eebcv6sWIScF
2WMIv4Ox9bbRi1yuAscm2Uijpn6JuFl2R7c5DX7txnbtBlu/JSu7jRBgt6GhmO8W1Ew4aKxItcJa
PGWg7L3GPu6vmwPN1pgDeRulfsQ5SaB/G6ZJyS8PWPT12LX8kT5WS8tXPFZ4Vipl2CZZPgHbpQcx
Y7sMjrgx+eJQfZVEpEUx7yYFjDoyJOJcFM0P95N65jhkzX1fy1cM1/MfhzOnGxKusDZQJWlJ7aJY
cHPPqNlc8gws+dO0zGL9jJR1eXP5MvoWSJmnp2ldiD9MfRyxZ0fTl+3zcqPqBmXchE+8VkxuuBlg
FSAwP+kb0rU2GCKQsH022Uxt2aWqJUm9ajDQVmDMNYyO8STmnhTqWeVBCPjmwbiLapEPJrDkgwdK
YVVi6rE8lwJ6t83Jl6COS1efpvAmJ/O8DCREzV7P2DD4THSIn5QQ53B5jDL9Q+lbthU+/ABFGC7f
Cg/iGCwIh01sTWtoVQ6QfIrelvMW0AGH3lx5SujAybe2/G4xgtFf0QcN0svnxfcpF6Xw+Hm663la
oWUHmISJyufzqX6a4ITDY9QEK9sx2nn+IFGpq511166RTYfb4PAIOdl9CTWl56xXPctJ7q0ZToIR
I+qaII7QMteOgzHLdp992EYweWRGTdLq1xfMHjnwVVefSyaYeTRbtf3VjhCOuRlkcXITv+xiVlwQ
lUWG3EcaEVZP30tui13k5FYXI5/JFs3nHCfP4fiY0m+GDccdPHn4wAvq0IuNQxPKN+ZmUsNVRjYq
g1H79nNM57z8rvYF+KJb+VVfRcPKgQkJsF/xHkJOALixsv61UMO9szhmsAPVO/Fq+8zWYpsrrF+k
IyHDgoh1RjHFxpo8qA8Gz5zNQJq25aqyoEZ6ut5hGujQr1Y+fWNbFv9nkMak8qM3IEkuvQmdFTMS
8lP4ade0a+qvHd+glsawGaQG5uRgw8FddH1cpUwZHvmzy2I6Vpfs4deS3pSXHjL31M7+6UoNu9mC
4reK1SEl3CSeWHQGCD6xfYPTa3jAdjtdvRdNkkZodZOAiXpTLcuIzgfun/Qz0uN/9E0HBWAiPs9+
+2Abj4AfB6N5RpK6fapOzOlfORxE+nnXZfASf03zPinO5v0cSgdrennlDzbg1YuHHHZSqmeQMCwl
ib7eK35JeaqDOKTqrmCIuSySkaoX7a0IYSS/M91GYRQlw/j57uP/pItCHLUzBG9oFUYLehsr0f//
c5D5Pargx3BhaHSydhGWOY8ZnsWJ8Ks0i+yoG/ZIfH6RXelzTLeWAJZSFg3cMSgVyPA+OQajT7+L
G60pf6/ceB7q2Lfi7NCYv8l0e65hyHA0RR5ctdMlaRpFuvHsVkSGr7sHvL7wbx/yzljJZ1YDEChC
IilVTh8SRhLo03NZUnHi9G24rPdXIDGHL+uxSzZSC0IdrLCioXCAWaU+CbEJmfGs9uwKnvae/ohW
J3BuwuEO0xSX67PtGSkCXCSxl2333t6udcvJTbgjHox83l3rs5uXhJ1n4NBUuo0+qw0TW7EDmSbz
tN3bEVBQoBRpPxCvM/mdFG8jrevZIcKc93lD1vhNtdohHhIp8r4smyqYrIvQSDJ6iqFyNv68zTCE
024hODknnUbpDgWb111oiXt7c2lZ6lQ0f64km8YZUCDZ6vEiGPAbijf17ETLv5g7159GzD6RpG8i
6mhNLYgl5wMfqN0rcSAF0L+RscpC5sSawvDRR7UJYN/6omdy3uYj38ey2E9R2MJP3UgNn3nW7MwN
8LGQ2lPHajPJd6QR9/xSNXbVpoivIhBD4f97Koda34mk9+FSOhI3fJfKGoZTWMOFiJ6eoMoPTEfy
rE3vFrtR4PySOHLoYlzdFyh55Cmt+AKyOZ3bcf0RMGRFvVSN+zRBjVed5xNxFsQfDfq27i/0KKVH
ia1ELGkGI8ZL0mgjrPpWQswDxjEO8qqoLSQLdpyYvSiSOUsTGoleBhhnFDwxRUeY482SJVcVyaQW
WPjBr3RusJk3f9Vs7wPh+NdUUejJyXrHuYoHbbjajvtSozzFea62cK3x5qvL4JCbSKREVZ2xEIKb
prrLt6Fiq5Mbs7nusNfWBB+pALNNpMglsp9Ipt6Iv4iVXFrs6tpqpyDQCaZfhpAW705t+YAe/Ap1
92/rfwVwo6JuQOmjhAhg1TPufG+CBIO3EKfMWtFuN6Ug3pYk+FIeAml6OntFh5j9v3F2Vqgx3NNZ
EcAflAjpwIxUMU0n3+q2r2giO/56bM8TCEwgQlI8+qoK/VcLmlu8AttTZprurIXtw6LLDuj2GxzF
cx5eo81lWD0dKKiMRdLSzcEJTgwRUNEzGLB313AiC6l9fnWakJ59H0LuPjLwrMnYDwiiKjVvaE+C
SrBCkqZXu3264GXV0nD1vDnI7/JtA4dFVbY2+hGTwQWv2sY02lomYiRgw5+x2gH+QN/SHnv1YIJt
6fsFyMFd/TL/55fXKDHVxhquW8dt+wLqCp6dz3hAyB2iqRNggWLh/Wcl5cuAr1wNRRXlNtEIGVnv
1jweIIhnfyj8dWI6UMSj2I33f1ZpXM42h+k/5d+PxrGBYWGvu2J72sKYZVZb6dmX7hsXEI20HMAq
MM5CYqmKEwwtbIM6p3R+8vU88WPtQc5BNNZ07LEZZsKaoQ4qm05Nz4p2qCAxQ2Nw8JEPj9sWeAXf
oUAAFFHhH34HtFQ3NwpAZx9z6AuTdQKclw8rFUmZMAjTd/8aF1JDRK+DlXCSqaGHVWRWqckHylBM
JowxRezcH5CNWVOQR61dKVU5UydkNynQ/1c3Q6N4rFwj2Q+ZRMr4cIWu9jgzlVRxRq2L1CdGlSUT
XDSLOML7NJ3PJD6LllmY1r5J6PBlxfzNUnHE7srYdRJKOJU5zsnNxZkDmyadPvegR+8TBwZCUNL/
Qdu4qxE3yAMOaLTNoXNmNwM3vbp/fOUtVd/PW1YqVfQ/PR/IoJraLcU8A3O8DVPPY/Ko4W6SDP3x
WOkbrm1BqUTSUM/87LnyRiE4BMzXwrwnByQWRFiXbNVrTUXdA32JJy8ZJvdI6X2N2R/6c45lY8xf
KCviXNLO6/9AnkarrmVxvuX1sOdRwzt3zu644dsI3TIEp+Exhpphyd6hjEk+q/FlDzqBYOIGnx19
2AEjjh1U1T2tGy1+7RQwVwVTfAgEaRufPrfFrolLAOPxDplZvaP42Ijt8v8T/6Jzlmlt7EVl0a9i
SKFqL0uzLWASx/mY8SXsrCNyx+9MXYfTEU3emu1rVyVdGqLX5JEiqzq4/q+DOhV03W5OK4efmTDw
2gSu6vsiduG13tgRP7X/AKckp3VRL+m0n40fQ+MWwoAqnzEKJ41oD+/yvnQ6o2C9xzZ5gYCEi1v9
+LuVO/oFbJVMgydHKGR66025j54WtuP0Hj5t5q5vgYPYMYApCOnYATra20n1Gsw4hhIRNhH2RUNI
YiW6uR3cEADz1Ig8xMxdWcvZONpUt7KpsVgcM7NBBMf19ovQXbdvQ9l7HMiK5G79PIvMKV1OJhbM
kZBy+S8gKx+aiYPw6VTWbrZJxdBxi+gfGTZnR7PJMdHJDxXAaF2MGvyoYEQHzFtRnIcnn0qYCNvi
LDz5v2Ypx0S8tKYrxdPn8+02zP+sa0L/DHjMi49UQgb4oododTWcyul+qYE2UQ/ZQ3lHnIPm6P5r
kvSFAzEQJnEnZYLVBqZi0wRFhWK5fLfWmAEnAlePccQNwKzc7Q/cR9BsxrQSQkYAyndll0Tg1ROv
8yQXQMbshwZbK6ph1V7zsTcVW4r2AownAkoKsuQoDpV0Qj+6WVRAgotATQpvbshuCfbW+bdP9y9c
2UCgBVYN2SyYsQsw1zYAUqFan+WI5Oh5vp3k9YB0zuVvz1glkEF3ur944WyXA8nf8F2WNGPVExpz
By5Qvd6gOUzylSgXgI9weJoMDexPS/5hY7XIu0AgpAt31ITI0WUOYUPNuRBciKWgjwCYQF7ojI56
pXITa+LQGk5fjij6C8CROedv73/1aB5Lg3R84yh3Z4c1kKQuSzL/j2Z2e9txNidoVTmVKU3RR9i3
pPFVcNBRkD9S0qD710EROIoAC8PRMpZbbIYgB7fcj5reV1HP/TsRKGjiTc+MIlE+l4MlpSYz0frd
0jfz+LdwE4/kcjOaHkMKl8PTALqQ4Zc4H43kCZYr9NKjblmGsxXI8QXRIgcduGmpR7739XTS5Cg7
Lov140yck73HIg2PUSnMxVxE26tx01L9/3DXU6MsPWpdfIh56x9WAG0lDVtDU3Fj87vicBd5sCAR
EJs6E4vVd5dVcL6cMOZ1wAkaq1rqN15AUAl9D/zbl16qK8FmHif7TnBsdW52yHKKVUzd09dF7rOB
fE401PRAJ8SCTePfW2ruJTvI228uDeJmg4q5BDuDcZOefLMVrSI7vfPMMdCCE/RULiD0CEyY1Tqk
/jFXoGpAvGG4A0iGWVQFaeysVxjz8VgnDKBmBp+cIH7UWI+2fBWTs41U3PTOa7hGWyXv6qJE3Gdl
cblgFk95UQyY280cwoggBDoGA8yMalC1fZfZ3UnKldMgUfAyp4H/D1Lmh6099AwdEJTc9IJPpLHw
Xd//CMpUwxaBh4Nh0XdiFCa0bEAnyO9/215CEbmqjFn4QQSvRxv6j3PP9zljxmjoSX2KvHEnsbQS
h0Lw6DQB8SmT4VrM/Cvu9ByXsdzfT8nU92y0SBzRP4NkRmAsbZiS9FfqGtP9uKINXr6lejgicVzV
sjhd3KbmS3bkG2UuYhLVVb8auPfkV0jYvi+Af2r0bpXGnFgCE1fpPbJSicdZIFH2l1/C/hqrdPed
eoFpoQvgyl+gEXyz8/4yPqw9/jA3iw8qAx9Ttz5sSuTzKJUmYkedBMKkgsOxabY+Bxiy/3LqV3Dy
+RwmLyNfzZdA2TTK6nZPWPwfySSui65emTqQxU2ZXLWjyvWwv953HJHTMdQwdY3B0HBaWtBhJNsT
moHpnbtj9yHvrGLJiEfpU5Da2N9F0tER99tf63pZsi+MGpM4aFaWp+hAfq8SVxdoiPzn36+WsXX5
362CM9hBOzelKwTWfuGYxM42EJ/++y91BzI2+YvofNFhbaxFR+8TRMBNddrAMr6pPAYy6ysTaE/Y
gntzocin14Bau/PThmum6tJq7XwMerIZ5IidH6lDysGSy0hbIRzl/A1Ka1oaMYUBgR4R4QbUAVpl
05qWCl2Cb7I5GzBmyvIaQi0G0n+wad4aqleAXtPSgvQEX9cYXOjvMNdwQXYNkqQo9oplExqih9gR
iRPTusBNhXBL4GLbVFGfHbLFDWHItMan57nJHqAqfbNpEER7G5w9KUrryBsdqeLeXAWg8e9ut7pC
+jGwI/UjmCSIaEuWAUzOpRjX1JTWhbX3IAR1fDgqP4bx2XBuc0M1RLkq9M6hQIdkVce7YzdOMJ5s
TFg9tQBmxuvX6WzeYzSZtS8u+DQd3cYhP9zQHVzsjEJ5o/kfDhDLwg9cF+tJsHEA+rbr8hg9HTVF
LS7gTTBM0hWGbQYiZQWdWVN4dCXWJBVhvwnMXwHiCybbyxIz5d1+kWpF1GxLAf8+iBSIO641IRtK
d0Ddikeuxt2sjqJLUhRZzge4AkkVNhzxvAB78VNCnn4HIuIkkw2yQt8xbxHnEXDNZLgx9XywxJkE
p5wEPhnlnEywpHDUEwzd7a/ATHcpIVmmRRzxJC+vYoCWg6IMV2dJZqu9w8BWMwHhAMjEiYh/IGI6
Sw466tVWWT0KcE9RD3NJW/j5G0AEODwYschPPlcaFY5RZeN/RFbQuAU125gN54YyESnNZhU05jph
mpUOSfDYsCiUdm7+W+veKZX8QiOPzoR4HcETkFxAViikpF1yDJ5zUOoarzenayMSgIHgnFvAAi3w
I6XJtH6sv4JLsdaXCmjbxUiXmcbstWqG9sddqrPjRLaV4YBU0OAA7jcJX2LsxVlNvjN0IYMTymPT
GO5fq7bYEe20gt9v75R/WGhO6/D2rxRRs1kuixzusadsuAGcRFcczX/a0LdJPrExcdAxbabJ4F+A
SHPX/9TzvtHKzR+7drxus8QutM9KFEzgkQNPs29YmtjP7rLcSXHwSPcuB2Gcz4amOToHeA7kagSH
85rM+1Yhnz9cKjEIsVuximNi+Z1ZcF7cRvTbVocZGIIWniO5e21JyE2ClO/XTuqNNeyGyrCCDpsa
m1WashyVT/HhaF2pcEAH/Z3PwCB3QQ8U7Dih2KjbAPV7/Fr56KgEjDp5CUJL698sNW4SBW9VUd7A
8NuotkkFuSQ2vJCupJmqTpmNvixDjPM2o6NY/hTtTole5W4T21UneVOcIXa15qt7oDG29SNUDdIT
H/vNlPU/WQWe5QJrtI7wTBekPSsy4wFC+sMMxRVrCJtuuEZp/Y7id36+UyBw3Djd0Ez9K7Xp5m7S
khXqy5c1mwdJIcx2c0+xmojAeN8dIvh+SwL5pL+1JeJMrj9wBdWmScOComE+ZsLLYOQzyvCj6leK
kc+u2HGdM4kZxSje4Xc5Bq16ewVuW63O6NcdYtwGvGbhjvNoNMKJ6A+EiI2ZdC/mqtCaEXb4089g
a07VnTfbde6Tka+mlY1Zji5AMTjYGK3fJ3JWa0ao/AIWXdEC2LbcMJQwwIyNcIRpFsrRu8Z5bp5F
ePyF8ll7DtlYDZfCMmoKbNFR1EHskrz4x+P9eq7zhe9U43JsP6bmLM48MhqXpXGJEq/Gk/xVfFpw
sW7fQUgPtK30x/M3gV1PlSwh1HZ4eYvPoxVqeXNSjis5xU81hc5PoYsgC9cHw3M87VY6mrbU+lpL
eThax1IPdjTaLwdSPxblY0Nmr0R54N/aLXIXfI/VK26E7gvcrtVJXG5lgqaJXkG4+6DyFuM/vzgO
S6CSQAvD7Z4THcM/2iJO1XS1nR7BAGOWUpTeMNcNBz6gXzrRuTHfut6TQtEo4CiJfgTYEkJf+4SZ
XPVO5L2vTb8KRj85t0vhJSRQ1y/9f6EHJE8f//gOkAkNKdqzya10TA1mTcBuZPRCseEKNmNn9KtD
/7RbJ+Vj57gm6srSNAo0D9RayjGzHtDKpRgA7OdQCZmAJ8NmZRnddaEy3iFFuhxGoYqMgV8Fnp+d
695g5H8Br/iJqwEcwz2Rn3YuVQpSSNq+ukV7/IeiG2JlbID84KD/toK9MsIoIlrhVlqpEEazFgg+
GOOLDsImY4GGbWtwYR/YdisfuWlZWsEus66Ssa6LxIX4+nU5pyMSNx4y/rU/OH4ePcbRQlhu+Leq
ikPYK2/wTRlkGofc27McGZ4SQZuuMK7/5HyzFv1zOdxVgr0w0tDWDpmdrmoe6IKTikmfaXKU038D
JIN7jsA2K61xyLz+PPfPeMaubNauU5amhUsfOsFMB3fxyyFIjku85PxUYpFZxYVSw7kdMehiDCAC
26ylRdPZTFvxwlka0vMajoLt8QWwUgjFVagZBVCRsRDLElErWP8fL/40VjLR347VyX4gXBEKGrA0
GXlTon4aGKkelfhoINbbnbxjCUgYNDetLW+XnH37ZO3fkFFyFYVCvW8Dgq+pdWa7uZNjZl7QmRFu
yOJppEefZfRT0zMoE5pBjvMcU3H8ZozozQukMbt7EKIYbq9S8K3SI/JRqDlM62e3W+IAJ4AC5p/0
l9uSgGOM9Qa1lqdDtsveUAzYGFFnj/2dqMZMCQLPfJg/OuVNTS6vu/KzpBiBsllX+rQfRH7df/5S
Q6Q1hgr0uus3z383NcQCgveQ0Cx4n9nn8m0JhMzBFMgc5T6Dr/Hi+xNBFaKqRonSJvTsRxaSTXvr
CY0lPjbPufxmt4qBuIIb2ZWy5fPwg55ocCg7gHfN/pofUQ5IU807w6ZwdSCWgN4IGlhZ36g2+7Hu
1am60KZqT86RThfC/zWEkL0pZKMnBy/usLH8asP+M8OOFnZTz/dF3yvWqy98yju3Qgkz4eHbazYZ
hCIFTwaQdWXi5oG8Ud2JeuHcQh0iOeJrFzRGt/kKYsjgCd+8Cxr85Xd/+lA3fYasDzsO15oN3c2X
HAdUvlO865x7cqyys0hWdWrquA30MdfA7OGsSY43FNtjG7JOPKYUoHWp7NQrVMWKvKnH3BaNnNka
AspZj/8ENTIA3ZdrF0dh0M4p+BT1PyZqeLINS7HLff3cJDyqsU8aT0gdfzNYGobDFby1Pf8FDvhj
StmLDBYI38I7319yN8DLhCjIIMK8RcBURCDUK+0TVJXgtRb1gA/3dbJXKG3X6uyqc9LAfFES1pQj
begymDYCVyI+BF83yRKp5Yypj7YkCNtSfIrwLPH5HzWmkFMd8MqKaXICJUybW89UfYbWCbxzrk1D
k3JdRdV2VtDH/BSQpYu2nGFEQjqRoUu/7ufApgk1N5MW+eS1Ob284LZJuoVoVclnF4UW4d+daqeY
yi5bQl7cIi5ZKg+MFR2xy/lwe2PgEcMSxMRp8p54T1xyeVzMzP5iFT4/NTufAFFvjbXkpasgMvyF
PXyvBPPtiDwLCTNfx6ljyHQATN7NobsK8BRg7zwSFUb8aYzyAGRA3l+VXEgwUC/I5xnw/N9X7/0s
inqTKw+oapH1tR9t/ON+8ESmFIAAdUAZ1Am9Lj2xuHKOCG22bqOKnhKk71I5FzF9Y/2kgI28/9J0
k+w9V8wQm8MceVSVQPLXyrV75aOI51oAH+cI7BNK3ELPGWzXbsZhSeQFWIBdJCNraaOsVZd9bdPS
5HLkjODmnZ0D+V0rf85R3KdlZdDWiLau/vOXokLxrX+LfBvwI7dyzMgE4Kh19dZfLEFobIKvrlUq
AzEm1yaiJOL2eQJFftAzuVHNRimaLMpNSIQ9XLtxxzUKYtYFpFUp95JD6uDuno9Q4iA5nUZYi6AF
Li5txbrIPmrVihyxhwyQeNRA3PnO5fwM92ywdBhiQ/1OmxJ5XA3lxMvcIqvgVSuv9Xq1Qlg5O2WC
rY5hqVzO6EVoLiu9ZMtni3H9x6wZzVK8Y4pzzwVlkpALt9LYtfzsoWJgZEAKoQzs+oUYtXSKwyYf
MrMQ8TStpBSWOlWa9f5ONNEOXLPjdKvPeMhxG7Nr2AhsG8/m18E1LcVebbj7dQPUeR1BaniqSf9k
uXQZvg1uTeXpEJopGr3nVE5rYdsyFkY+eQMpu2uRUvTx9wIvimfvlnG24sgfL0LsjVFYwxvARbHC
QlRHudKFECdixKiJYBDq4wnAaWNjBrf1p4CmZI6wZ2w6wQC2w71bnPHD/gM1PJyxG0EVy5L6Keci
aJ4bav4S7+KuRVhlHanzvC8wKy/P6drUev4aUSJVb23u+uMThnrFzHonD1qmh5/d2T/uRta0hRmj
BqyTziZYncYwg0Qkg/vxKaM6t2pQVVcVkKqCvTuJJjV+OLfDVgw0doh+S+JD3O3eeUPLudRM+LHY
82hGDH1WQYcHylAZq4XwtCsZrI+Vhvek6YyJYeBZF2MzpkBpBto66OXyGmSF+g8E8vumF3TIQpq1
z1JdVCffB7xv6+s0DkMGpNyIB7ZUauhg90NlO+AxXKq0aj18PZ+l6As5Ci4RsYhFEYR4Aj/IEkCX
XllIejtrlPVEVYdd8WGkHCsJqj/99Q5TdBzBfOoHuJJT+kQuU7MJXiXKZSQtIOinG0HMT3jNkF76
Ki2DRq1BfT6wyv6dw9ix6locVlAjDYtVsG3w9kWSYCkPzUTN2+EpgnYIXSbz1zMQafCpcLQPNGm5
01MWP4PHIDSoT/nrG1KFAP/VqHG6CmMvUDHmjLbf7WHRzEkcbilt94KRuuDEOJVvhbWa0QCvDVd5
CLn5YX4G/pgxNt55FRBdoQEC+mUqqAjyswSOjKV83a3F3EFEtCH9dfqGl4XXGL9et8CJPPwLpHmU
7HFZUtHnodaRL90PmvEj33UuJD3BsWxoag+sjI8K6546DGklvF/Ittj6zLdAyb/1zlbW6gRE/PfD
kAXyQFFVJqFuIW1OMDUX7ncpxkC0UZecmB8P255ApV2HDOwDN0UIWxZ7RvYczwEFtaKHx6/kcn0M
0o6u4ZBLDSG9TBfq+E8YsNOA1MFrc0fn6RLhhj+29o4n7ekxpR2nDaOe8Z9F+Vn0aehz2ayFJRiR
A01s2asyXzDz7OuvDHV6pVMjzKOs5w9mrYz1slb8VXcSJ9eZEBLzxLnYcLS1EBgfe3hhlloyFyBL
gyJEhd53qZFbubN+OY6dcL/n7b8ZTWUsTjppxgUtIpEWT2itcT7k7zuM0gqVbvZ6lHkFuGivFRqO
R0awailzbSv916RUa5JEETbSGQ96I+Xy5swu3T0WIrFAZGVeneHvnVMsWbkk+HbARLwZskplv1DZ
Me41AJCx1P73JMwYJUUiJa3BU6EGqUe6PJhJ6qXbURijCFy3fl5fryef1UtE0sVbeH2d4AJACaTL
qvOiweG/QCeLmuL9zKixb2YNGcfU8cq0nYhJafd1cYd6v/8vra/rd+Q3zV+CgxBcVtyK7b7ePnsL
cv0sm/PRNdeK3UmqN7P5h+MzwClSRrInASHRmYlGr3lbMDrynRuiPsTN7YEp3kOVMK8oDrU6xipv
eUSu9N9/zc5MNvWhy2ITm/jsYqm37aj+bat+xGz3c7QidFALlddeVoHTnKARgT/Lrq6Z/a9mJsml
W66XoW0uJyCUXKNxB3+F7qfjr7tMamPFmjmcPQzxChe+Om5end2gOR01y1Y0MFE76AJbRj0qeZPJ
eikda3UgocDVS0ZNMZBuEcxXb+RQsTzsP0U5unZXk29F057I169v87KKNWpj/lTzRRFAYOXwgTVm
2VpDsHZFsk8qZ5D977FbsHxcQu7S4kkplKGiyOZw7kwc+j4c3IaAP43UrdpDNNIqYJtV90kQzEGL
u3P8zMzf/Lbk3O+HJ9u6gp2qgeOfxOpEqhW2+lrk5OvgWbf1jcfgGPxfqUtVWX7ka6pzsvIzYORs
BEjB0QNVvyhEdbbYJxt1WEbc69QPu0RTbGr6U9hAmej3R0TeZiFAfslgjs98By5q7TkKO+0MSrWM
M75HrUNJa8msE900FJkqTV1e9iGAWcJJl9IsIwMb78rvSdeuDvEBRezY9sNaZGZVQ4s1lg1I8SqA
ctsN9/zewbMC37gxbkFAN6OPJRdGAKsMNLOf6Fkg+ZgA9G/xN8gDNbvPYCMYRoK+avrhAmbdOV7N
RklLdwjNAH7UtEDoUbrmJxjpiJKmI0WnahDRz8oq2gPrBAwPCTWo1u0XBE4SyOHKJO817vfWsKGe
kaHBRhwKWQDjQ0AqC63hato2fB8kp9PtzY3+hq5aqRLz1cKMhs3ZoEfpmY/91LJR7AhDrJ1R600E
l13sYEyYheFusFc+SJ5ipfzDwvuyUIH/ssF1gcVcOpTS264EU0UnDOfecnQTIt0Mo4Mo91n0sNW4
HE2M/Um+Ig9L+pSt56yHgRc/ZeZQ6yNgV82hDIbwGhz9jASNjNaPJpqWdzKRt/JRrSxqSDv6SVOL
Dj4oWq3cGcgvQmtR1y5Bzsh0ArmjWK9xMWASWGlaSQQjrJQs1oMJi0H/AhOo0JIa+yH3HaPgqGbC
U98agLX8dJ07cZ+YubxzrCqyl1+qXak6bSJ0ABxvDNlsBOhUkLhDQAvIGIXtLeo4oU13KpvurzpE
iN60GQeMQpONuCOwr7OrWG8aRMhg/F3DHI78yHkYMJsFPZ/QlfvCLYV7JLizlNGJIFRhgGkj/LpF
3CM3Dv6HX6FE76wF+TJkKc1ZwLME1otOA/+lYud68Wa6OxonsF8oJDu+PEZ5YLaq0O0TApuZq9js
ipbbSCszLVt9xu2yWZ4K9kHUBxxBn9Xhb6thV38o5V5OTP7VOY6Bt40Xb1sbjaLSct9IJH7Qgket
h0QxDm+T15Ab82gkEu1ykOt3V9eS7/Cc2o0skt2h4RljZU76jxLG/3A2dAZdVGiCzh6HmBXOx0RI
FiofqXNF7bOR/FcaaichPuRUQ4BxY8OLklYiYpPQe1M2twnqKR4MHvBsh5kRe1O5KSiUBBv0AX4N
bGIOPYx9/vK+7Y51q696oYF5v36BF5uCh81CN+nW/VllhuZGtQINMeBGP4kKZ951e/vthmcDp/2j
IGAYfZcbaPHFAjA9lRL3ORyF6QkwlYSEiEwms3fdmZS19ZBRneBK0C6YsbolIm5jDOlgfF55Ut+S
HiyOb0IRpV0jeASJy2YKQdYL76iCbWAAf38cTmlFu1ktZ6njI7eMT08d+QrXuq3Susfa9WzcsfVQ
nX8w32+zdV4NTTpuX33wEsQ1tPYofMZv91cCX4R/1CvKjxCmq95gsITyH3DMe9wOMU54ABNlrJb0
+3H1oBZfVC+u9afFP5Z3pAor1ctPgb+Vng8zBcwYwvh6/5KqROMbsvmlhkyhGJWaQbyqM72Qfys1
HflSWrUcoXygiYEjpa0ZPIgDFJxhQtA8TpCcVxfIqSR0qX58FFQaNmYxjAym6BhFsWCUzfNiehDy
jsCwXNKO6mUkv8k8oBWrB0lxdwRydTZ2QMFUMJYdVwaDfuKEeoOiZ80SkkgYMyzZ6M4jSf8Q3r2e
7kl7rfB4tpQxVf4DfQJhSbWMF9U5qXnaz1nCilZv1PhJo4jpeUHrqDM1XN3w0o+pXk9dfqkIUmOq
ih1EVkdzfVdwmiygPKko5dQkLlPBhczzD+X4izNLZtqgsVFaTJXaA738UaN/o1zJj4JKmzLLsnUm
g9qTgcIuPT/8N7B81dMnJx1Uy/fJgYnpSMriNbQqDDISRF8+czHPmt+0fKoFMZS+EkxCY5ux7zm5
Bnte6qwSYW+jdXhwJwwWuBZgdJv+5Q2yVIYIfCg8x1Jv9y76MUz0xffCKgwDYK63ZRX4UuxRmK7M
eApUTZxLcRuN/xZrivM9ZCJCfYZD2UAs25nXkTGEfUjnRwlPaKSJLtNNigmZaZ8ETxkjduw0RleA
Nwlq6RbRAjdUgbKdXzBFCRYwQDkul4p+JDx1ZDh6YJTo1/ZCx+8OeEBs2ZIcS7kDrul30UBbMZ/Z
/UkJC1/+vRFcVpdoCkK1yXoyV5rr2JZQ5fGxBO6t6uTaGi8W1tJV/JMcVaJpVNsrK96NFzfRAZSc
AAQ+y4k6lU+PFWVU2p6BLdq6aaIWQsaRBkc8JTdCIJ/mItMHw5YdMbQmkm6GuEOCNtO7EomcD1qL
/aucU2611sKPVjeesGZ2/Fh/gULaMj/wZanERyGE2I7tVQUp9+ub8eRLWqWb1Ev5hkJKtAUtg4l1
09RuK5QeqghLfZrIH3BeNCZuluZ9YXFlAuXTdoFUKUY1elAyRYLnJOGbyMxwPaTU4/zfUoW1m99/
KBhS//1O8LnxPokpp/sBwaTrBIZhsfGQpIj680rl4/nCXrmskQjYHEk7wNvpjKwf0ACjgYBZvREi
kwLnpQIjmwbzglZxUrun0ASu/3Jb+99H/qUCaAWhUCpj6Tuaos8BMVwDv5jTvvbM632GIs8XFLjL
f2K4aTcvDyzt/6pJKIeZGSrPvrS+sVVoy55gSZPtP6AiddIQhNOdpbMYDdyoGp8WrjRU8O7sZcUy
mhDT6GIxlNffPT8mSQxkzDJDyCrlMq0LKvlmQPC39mFqE2imMWNpW1oRhB5T+pxECbvcbMMKwjI9
D12Ge6ccY98hQ80c+Vs4lTfwHPG1O3fVv5cH3M1+u8QXzu9TnqMuqVqaW18vpnkG4sa98jDB8NV4
i5NnN9GY62mXytzhzV4K7WtrTeeIySUsXQ1JsHVdR0XrJQIg7kV57BbThMjrgPsbajyEckdajDdg
wdt/7ILbpafJtRBKfhDiVeAptE8WY0r0fYe6aC8e6sZTP97tSZyn7uSIJpOhYi1J1fGjzkFYeGYN
h7upYwbVNBfDheReL4uA8V/GKCPWvpRlOtJSkvW+Y7Znj73OTAEOSsJllljfPJ4ftLGLLbbn6ICA
1iSeQ5KHz+SGIinUbqCE25ESmjr3x6dmet2eLg4ViGX6Lt0cFzaNWSQcAS2xUMidCUZWCZ8Aw50c
3WXDJVbCDnja8MiJWVofgwc/DcKjkzddlyGMxj4naItOfd3W4LRl/0DmYf17GK3ZfLd0B0GwfROv
BlMJ9zvaj5cm1EjCBR+vixQPqj7KIbabWkHKtZxVazOmFNL5lc3HoEKXeJPJVLjEVaOb48t/r0Pv
o5TMNQNK/Tqj1AdE7HU6PFFmPgzcRz1NT8HwbGZ54Y/WUkJneX+phFiPFjMJDA7NrdRSQbG/bCWJ
RAN0vAW2UVq1g2oKLxP+s43QUwd2rEQkav5wrvs3ZEYFRYq6U5OPUg17R4QEWr0rR4p6FLEIoZMG
++fcHNRJNc8vG4ABDjKaaMyXtKBlfIyiNlKXPlOAMWYAB/YJnQXC8EOnIEavyfTPNPwSvN+OvLeJ
k+LPJpvIcOp8SHiRKy43/L5wX1bxz5EIZdpM+QW/+ZhUsx7Pz09cFClv5ZtbQec339iAEv4RZ8ck
pC9HChDZixTOqbShqUZu3P3PUFD8ZbgrN2zMDmUH/z52kUNKJr9Z3ZXEiRybSYoB5CezPeAAhYKP
7YsU2nZsL8aOnzHNlHnQsAP+40XVQ1xClg/8t/MRiLozsqY6B4sFbSkZGdog3qW+x+bpnWfZYS5P
pjdcDWf6Z3J5h8ygOY8TZel82XzZPsyROgBnESJ4cZ1R5jNlWY/SBUsWsRpWHt+V4y+Yiyt5LfaK
ugH17oBauN3UjhYwTU/7DpSZA3etk1oJfpy4ZtI4ku7gM73/RCc4tOcJ1VwuqSa7cTtUk93qXYHE
riqeywOSIyU8PQGXJtuO04nlQhuq0wWKiOxEU1ddseGSCpWaAr14z/JAprl4TlWAuJbHgviOXVXy
ryWZfuUAi6zzQDjoc5UfXJoP+/LMCGw07Xwl2VYmmIQAhEkgrglwYIWfiQJdfP5wABunjrzJBDRj
oQFkamEnzAZQOaT21+FmaISFl0JeATkLTvpjdl+3xKiocs3TtoR3OSS2ZPiLd8Ix9X6wq3803F6G
4mPl7WLv0Jak6V+QD/nav4LvAcQPLb6k8hUPfH8OKRUlzIatmxc3jLiMrYJ4RxkxrTWAPHQLxGmV
xFsxvErWeS5gNUeKDkrJAo3GWxzaQvru5JmPWZgBWox54H1ylUgaF2clEeSPhVxqzzoKtsiu/j/A
prYqLNSdxn2HsKbDmuNXCXlqBQRIaCl8Lh95Goialds0OG476c0OKg/LhoornLguJxfBQvSTMVAy
RhenkSKe7nUEx9Enwf4jSjhoYIbTCNwSrAwMlDMZMeSSPERfccz/SkIxkS716gtaaOkBkXhhxt3Z
RL1LK5N1Y8F3ToSVmQHT7Iw5fa6hHKrX2UY+T98B2REixFDpsJfCg68df3BnOB+hP+uxzbQSjwHE
+mN4WcPnqPKm18Tlzez//+nUC2dj5z+ctn8/mvREs2Jj29W804VqwPXqSl7Bpo5CBxFc45bUQ8UY
Gg3cYNYRnsQO60JXRdhlOTgunw7rHow64yzE+hJ2n4ZpYtbLs7dyBdr7IfJFrkLE1AvLTc60vmgx
TBlZngkcCMqldMTz85iTHsfJ1Clj+5PFl59koKjMIr6HCvFhJpAmyMWkjISzgZOcIYUAf68Z+Yv7
mPJQD0FjXQr78E0BqS6YTdyWRNW/FtP9GtFyhQ9OTfoQreG2Pc4Shxd7Gb9vufO/mhvIxfSlFnb5
FkSSdowapXhN15ZGXdM9w9G4PbO3hZEWVd56SJGxzQ8ueuHHI1skOBj+jfkqOCz9zf552VyTQv15
aNGCuJWzfIJ/FFvnvzulaMPK4jsPCFEAvoaQd0qjKWJLjwuUtWUNteE4vtWrCt7GSeKuiWZZTe7X
9KoR9ZvNFa3XOXfvYhqsvH7QDwRyJJguLaRCNxTB88FhqY81sHTX4WVPBxFKmPD8eSOTY4Uu+Q7N
iYWIcBeLockw82B91u8OllazBC0wouTWJQL+THcT29g+pGHeF76oCbZV4YEJOmkuF5XZZ9ISRWB2
M2zsW9vDLFUPrDZ/yzEqxR644AGw7oL5hsyCILzMp1jnmlZJ7sOi03YImkTtjlj0k8/DTKye+ZX1
+dgyAdn0U/D6pA20FYoZsc/0SW4TlKNAgz/czcZlQwIRH9NWWEY3tZProIyFC2FfjymphWDpjyXm
LTXe4kcnCzYSu8Hg8mmlb5PA+gie8QS5coe+TummhbwxOFzCfNdpNX85J+SFJNmMIfNh0ogfsAtA
fWcMPA2pTsJO7mTbK7rwu6cWZMhi6AJxX1UWvhp+vWKZl4H4USRKAZuF2TkLAuPo5UpKHIVofNWu
exTuKWnHLk0V96wXbU6R1E1OCWHE/MxbqsU7ZPyqCLr3shih5u9lIdKEIP/nAeSm9VvyLiBc4OQ6
Eng/dLkfwPeZZbmOfxg1P3pEXpboaRGXt6Hogr7tZIlsxogfZoN2nkcEifWqr/DJxt4S4JvrHzJy
rRVotJ7Fi0CyNXUmgdIhBDh/xuuEQAM4ncSlkUq8SM1CkXwYHWoJI6KLy+1XTWPvEbKO1pDMqO0K
OKwSntioGgEmDwOBk4/DmxcGJ6eY6hXM6jCOX1z60fXrT2NobUk/RIomIsSdtp4uqI3F6ziEVvcB
Ismgylwlf+gZtbszp1a40rfpp8wKVanP4sSICf1qBljtZGCh+ditaAB3azncoE26O4RG84IkEcBs
QS4yjMyYK5iCa7XcQcgmOE5Ujt6HZJDa8aSgrc0YGTBiG+Zh7K2uMDnKL9j9lM8qCYpB11Db/oO0
ir3vXrOyD6ovqe4NOXj4ajAf3wvMUZ6yYIvfw9b/WBlbEAFS1iZjJ8YYz8NmlAMRictbhaeW7veC
8kEZPb6wJTsd/dZiqg07iZMEQERyboGuzC3+2yAGSqxrHGhvV2uX7NbMYKepAhIo7LJRihDICWbS
z53T/EST0XSmM02P03toADYt4sT10xRr5VqbyR8lLUyDVViNKeRuCnLZ8AIaBZo8Txeh7seKC5g/
yfv9uTDcKiJFRp8mEoGu3VLpaGKOdZ00r5XpUb9RT/eUZZR36UdXCTLsWh858hYtOr3iHiKBiNGf
rjHkpikw/DAo/U80e6rAp/MKavAnY3cgjal0yM5S7YijnluG9VxX9oVVy/vEqHXyN0xUek395aFU
QewO5G2rVsg3LBk85Q5WmBB6pDilA0VSYLHtrcD/LABnVwsiqjaOxkDvVhUWIhX3/v81yKkNVcjF
19w4dHI+Jc5nRWA2+es/v+QToBP4QrRZMKsf0sHZTjU63DvYXUVjoxQnRgxVbzU+TDS7hMKnl1o0
TSz47gmQM4esz1XeVQXS4QhukSgaOVb7IhM/zqfkAIgji8SALEgo3rW+MyVh4CXQlSdiETBBBlsi
cco39qYfZj2PmTktLwIo5w/6ca//3hPju15sobCNoSQFkRzOsuktpm1sZflDe5o38/NL1hcL5STD
1H7HohB+eIgMshyFLOLPL5fe3WjFJGuOCBwA3rFg5VeEs8427eJXP0k4BJgWgqvN0XWi4e3QBpxs
UrqA/9gJoUZk7YuJ23CfA5GrVrAweS/4iW+QtW8xwT4apbIPaAhwgqHFXTBtC6ad6KR38hoQmb4i
X6ULaUoQ1rlXvTkVH90KS53hFXKURQeNeuUDlz9NFnwMI4Ih8gPsYI6EFnp86/d2b/gvXJ09LU5p
VB0yFp0HUhMyux14RsprOUyh9t791zk+cV6cK9JPcL73CeGgbSTXWOf5Oo3OIoocbAf+yWCv03mU
9al1FTUI89RIv1Tfo6vPgbzs7Z0jA32ECsv5/BtJUle+Gli25ymA1dCkH3XMcxSnuviih6fdnoMr
nowDBsMX42mJue7u8/8tgn61SqyHdkPxE2VgmeIy/Km+rZdbGdEDpJcLsbweYr9nl0qH77NStG3N
E5flmDrgKWcJndb4ptPQUC0pKlqvZluz7xvUBvEVxQw+4jHzCeLsO//oPyIAc58QuRnSVDHyiwzi
EldEYCLKQrKy44cZIomLwMTgISK1V0bxJU7GO3bm++faOYYMCvFRYvp8KDcgwYYQGc7Wjin5TPzD
WUD3sm0FXLLS+3VsoIz0uBcCc5khEFmP9Z6aiW6M73npB2zPDD/+aTYlciCYwauYeKWBMNwyf5xU
dj4ko8lLop+1BN8VwFUI9x2ng+UJV+iYPpUEraD0f5lNLFrE+twWafvcovAL54QCIcr3ZHCOmItA
C7R3eOFer8Hjo2sStvihVUBmWQH6pBhT9QUY8jx+yzfzEjkeahjb2repQoqNHRRAtKghkGxGpQos
9a+C1H00WpjxIi+N6VgzgfCzVHI4P3hL6vpYwdr03iDx50uaTcZ0qR+lTem17+nrf1qG4Lpit3L+
IBk/8LqeCsTEqCu30Gq+NDMQGf8o/zTltrxy71AW+XO+RXMm1d81gZDSRJp4sFd65JrlmRMa8hhB
eq5FYTHoUZqkeV/bTE4Jmm0BU5yd/+8WdkFLMUoSczm9GZ7NfVR6m4dCZQVX5VG59cwFRXvrsV1s
E1Kwp9vkfnPUs7w10xBQhayUFLvFSpWx0/xVzfUEapFZFLq3SpH3cJ2j1F59WQWi1afg0M8xnJ3a
w73PMfIO1mvM7l6IEWX7UFGeCAdZ/aCm8t0V8pRyVSx2Q2U73D3WpM/ZN6TCf+DM59WKWTQj08ET
+0uXfd3aoTPJc8JJeb3bGEv6ZTvND2a0QBY/16UAD//SW3o6vqSGfwjS3yxytD0HRdjoAJGIhZmV
1B9fxClHRZGsWp9P7D2TDiwWWRAa1nbci0Cw3/pfE2ZILGqSDRH8ngeS1vLeGDztjexs7NeiqMMX
kXAELyou/Azo5q++zZbDGKWdvzN0vkoNAfrX3Tx37PkcplruGXr1+6jtjMCebLtCKQmt9HWssTN0
mj/zQ+9JfSF3kHJIe8iZlD+MZTlx2ZYU4o31yUtkJoqerFY0MJLaguAf7vjm5kMFdMLe0kbpx4o4
EJ9TSnCq6EOkMshB3X+k/MBL3wRYl+dno3CP4kA5err1zy7uSK2VaCG/YvDdEyt3z1ISAO0Eo4Sq
BV+K5JPHVOFkaUD/guxRECKpdaEu3UGKDmCa8TWH/L6tvu68Lap9EcXlG8LdpYP1ygE0BquEYoib
kpOq/Mek9k6Agyn2Kpo+utmHqz5MHVv5utk+BV5+o71q9s4JtTesgQzihsRudSrmqTgTKhnpnaGo
nwIUVPio8+N2ixBhZcSiWjYKNWqB+EjXt2zZRqp2L280Y2uPXxYpAxmaGiYculDbR55gd7H+Hgst
MEB0ZKZcmH5/rbzJ8Ou9hP7ZWYYOnvvfOXLrtPOoOCE4Lfj759+zdoPSsPkX3tXW1YHMV0bBeEmX
Y5GrpSIraG8T97AiJZT3XX4iRPTrOQ4sRcYPBQliLjfzv573MEB209lpmAlmDZB+yGJ8edg+Holb
sMOH7rFsnePAMBwLn3FDIOzuyWNUQ/ZWlKbQKOP9Z8XoMInoKwCvxGJTj0JH+dRI8iQldiTXBPbZ
2Ki8qq2u/OeGSZ0FB5VaRPD8RMB8luFRuagFxQp/2alG5+ey0WJG784ySzXsGTkLM6YBfJYmncF+
E+3H1hxsuJwi447TKOs+91pUCRBa5L5kggPBtbq39KrbNHPuwu3cAHY9mLI547f0D0DKIIXakTG0
ENl9nSxIEAkgQmTffGbeEocZASkJ2169VWETfiJL+cKwFGbhZ01mm1TWNreGn1MGmPZf/pBvDmVe
BuS3K57ol378KiaxsAFp3b7OMKf25ImLIugBF+Wn6pWHaL4KB3hvDMpegOKieRTxQY0IS7AQCV7s
8TUueEb/IXg4USYJuR1A4BeWefg2dxPXThqxJTfyuAaum0mWvxb/pM9finAbhgUKTTNFaLn+GetP
q0FANBXJBXtQKOsgSdhLg78+U2V/9A+pcqjfCSvkpW1ZjELuqE5qkNvsypt439b34bKCHGTP42OW
cwh+/FV8uRyDv9HFD7gm2EZJuJ3DNsM4CUtT2D5WMvQac70xXO+Z3ZgD09BShn1ljS5A/KKrOr74
HBVZdvlMvzZE6HqTNOlbkCzkDx6dDFHf5KEE1rWc9YHQ0HMx/PtHGlHOQQCW5BMZjshFKlUcnblR
TtfumR5o8tJMyuM/kZgbazO+xy8AuI4OmeqvbewmXEc/EEev/iXWDEzEetmOYZRfkOql+MDfDMO7
uBXcsSkjDU5BUkUM/zC8zALDH64HklZRcIpmnFE4FfWYWgHaG2I/E9KMfuCL1sTpVgcCRbQaPRtQ
abyuXorDvdmTSEZy8rIhlBmGlTmOzVrddeNNWcHJXK8cxgjJeBJ58bQIlDxIcv8M+OLB78VWUcH3
pLMzwOU1fB15jXgbA4c9MTgNY9uerBgvve9iaNqKqkcZT1O7lq2Z5VOU/jK0GVEfZUA9NxL9zu7t
Cbnv7TF1YWCWDyMEB6SBX9q/QZC+VP5Z9LHruSEWcnKM7SMmdP+IRzsZHQp1PBVyhgsQSvOA/DgT
Y0/g7G7+HqJJBrHwcGm5BjnlT+v5ihFoO4TVijYvm7QWkqWaykK60ejLYDP58wSsdlXYJ9azDmba
z3tLpNFiNEyBvhnokZYiUHE2WfOJSruHZJvcMYC8hs3Da13pNATilIgW53f/nydP5CvW080gbSvl
dTVA8fntEL0Sdg0ZPRotQN02CVkMZ5ycJL7z8WGrHGybjqnBEGXDVtoMNxjmuUJlw2qCYB3EySV0
CNWv/FvefflSYfDc0HZXkxN2U4hrGx3q+cKBB/XfwYr5O6DIXPghOW55HODVE89SWDSb+R6zJU04
VMBmWWFrRrw5MgP0KpkEwKDcSS8yU9L1qp7gO1LlaA18h+J8AZ6ctGRaNqVjYxha8UVC9cO/k/R2
9VtPo09jUhOKlobp3hmtJqaa7scEVPwm5eEhTmJfG+EXuuemO+B3H4eWlibM59OKkQfHeSml3Rki
WUqxzUvIVaEls7u8yn+gkunSSEl/AdoeBVOjibTxE3qgV8sbN2n2BTBlQaxZLxk7106RGEJUy1Cr
dDvAFfhky86K4K6S3Upn0A+6pZ1XMPz/Cz6S6kYh8jVg+xy6FjX+SXSKGWn2XjaC5PjPTTmOZXiK
/+y/Z4vfRQGIYhntmp6i9TsHeby0EAT5IJYismc4zeNlz5Bl5luV2RXnUM+w4ImQiA8mE0+X0U30
6svznjHyy60cagW1V0NWFVfG4B/rEpeAAtVoWmYdkFokgKddr2Y/7bSJYtP/YZFLvaZW7jWutPDA
rStF5FLWOdTFa4ptWwk0eVkSQZMLJmqslcNsebiSA+1XgSFCVq+D/rTzySn8RnZgI8d9mcuKfbpR
uLooPDcNcSXw6YvkXQNMqYWVGv8NSWKuikJguKhVLXv78MmmltpFt8Jm0OVDl1WQjznbj5qn7GjX
790rwAQOnvUirYjLK9AADVmokM3H7lbmLJmH6DZPCRVX6rX5FEfUXyhzDMF0+LYqMwenMlMmZMTR
dF8p0nRRNax0OpaoUUSGDYFqB6TIpvHbiBRC1WPGAXHbAaMbG1NyauuWmxMQGI7n5DtEf1WXoWOL
4D0lENwAs1J+qKTPeM0rqwtZMKdYUt9+IU9d5RSKj+YQzd7k634jYfUDvH9nIOF8L7ZqNZVy7AlG
24rJt8XRj2++l8Ye0VEvqpf/xN7bDm2R+wERzHDctGNUVoIqloKKc95N56f3zIbocZNvWdiuhPDW
ssgRE0DP8HMKhcAHc74kiWVhibA5RHqcOWRCHrImBY1uzt3tA2U13u71b5c3RwhfCQMWk7Sr/O4g
/bI7xh0W9wXqt1WhHemcw2CaCk14IXF58XiICphi7EuTWDFK20RXwrAMJjssiM2S08wXqzgEEY/Z
LLMPB8j5lcBe2anQhRFUMva6swhKSFOUw+FDzA77FCL+BNK3xkgaMtRq4mBvjaqZLTBOym9jbGqT
qAmAYvptfvd/rEDjeHJXNNsIjp4MMfA8QJEqVN4HxK04oiu+IZC0ei+8fXNqqQG6gf9Jqj+xjXbr
QO9D/59LReILZraAtfXRrMb8FyF2HfVzKP7i/oCJgOCq6oA66QuuolBJ10D5hRmKj3dyLtVq3J+Q
jOBsG5eDCqmdOO/b5i3Ax+KqZrdu6PEjbX0lWaQjDLH3A2uXcDTo7IJPAwBU7RJK80Oe4re74qgn
uqFtOxkvuua3wJsRT/uXzGcf+HM+sVDk96VIrUzFiayn1dJsIkA3L3fLZFu09DcQGQuvY60JGY64
WlwN0c5t3pRhwL26QmH6ZE1DTCLgeS976oOBjB2aqDtUxWg1dZESgXQ6Zlt80yf5SDcpWcdQOhR6
4Vh7KewZVY+BKZ1D26IQq2BNIuvyVcKEGUtkX9ZkPzfiv8sbHxbVp1nq78LWaJsn0BLqz13VWsS6
SnvazjjP5WwAg6ZUkA/7aGHVhuc8O3meFro7fSB58EkWt4B/iHFKwRy4pk4vBCZNND87lxBcNmw6
+28ulWYXDIOzcD2LfVvxj1iz2s8zSHGfisKiObskgm1ZPSqzpMZVWY6rNKiVbc+Pia38QKQlGdRt
IFGSRVQ3kObGyuy35QkjckheRJoQF+HpnApNtl9ea75oOkp37oOGd+erRR67QKD9QyLXaQuyauH+
0MpUVQEyOfiZFeaiBSXl3NuWDcWw3enzAR9oFoIc1DNdcBSlrfH9GKg44YEQmPeXasaQ3O0Tu1cE
q55/aB2tQH7P/MH7sorJjDU+gva8YheaS0aMvR8h7HyMjTsFQ43FWCd2IeageaD9vzTCH4PmXu7H
tk6WY4LTAVC2fNjz+F3BN/7bDlS6BN6ftE61BUA9Mrd8JGJCuSR9JKZZ0FMtjUuWjSVUjHEsm/35
0sW3v0ejw8HB0O4r3k8yF13g9scySq5Iah+kF5I7Bayyt/CqFCkTlp8KoXunDQLYozQGEwJvI2QM
2ERlIRI40dpvetauwrpoRL/8iOzFoLVfKy/lTVTQMX9htpHwn6FZMQHyKL10Ud1nmS7k6KOrqI0p
fSauOXd/TCQMbKmIANB0k6+/W6Axj/6rqdvPsqhWGMLpXlRK6+MI9FVZ47MirtmZamAnwBpQ2GA0
2RRF/pPTW7RElIhOjpGFvNxVhajFLAUVZIk7BL3w9e/Qis1UpM3uoEJitbHH/+2l+qpoQ9KNddyL
BHprAF3JJ6zmilvaQhTysMCLlX9PWtl6eS4Soui49utS9G0m0eqsMV/N9f23ThhKwrL4Spy+OURx
6k2kDbtfbUcIqbrvlhOB4wzCHR7CPOq9shESfQ0Xe3VxCwWuo+ycjZevUuGr/Ds0Vzkf+GHAz67n
LCa/c60bGUD8vxCZuH4+SlnscDn7jlRuPJVDfVJUrBqzLaYqrhqG555mNc7esZWTH1/yT+ejkFeh
SVLwd/9zn2ODFFKsrLFfOAW/nyp0N2AuHNpB4QIrah6kJpfVfLxeO1zyXSF/eiQT+rXhFTrKclLI
ZqY7rF9HSdbjKmVRnIO4EUblmcMIHVyW9KJXwjQcWG14A84BvMdy+u52HYqeC885DYGr2s8UaG44
IIq1w0A5y31e1KvcyS9zG5WjQMLPyQqQs81dPZF8uvts8fmdF0+K7EjayPZPvpPzPp1i5VOt7kJm
Mt4jZ5REDPR8zapIOy1vmuc6O6Vzdn45ylP4AsKo+wQIFFmW8MLPpBriKR1BofcVFelhP0+o7W5D
C286Je2gBnQuU2T8Zebsk7uq6CDxvbdMQWZSBhzqau6VbMx0aL55+jaQ9eEmWrCxvvhoWNU89OxI
OtgtjmicQkdp5Vt1U+t+2s5sbi2weszVcLJ8qBsxxoheAia6pyVCCIT5RzH4ztrkA0nRnb8nA/LW
vGd7yPGhAjuTbJKPsh6D4cJbx8gzVLJN1pcIjM6PBmiPYY9fgVa4m/pjMqYoezPV+IXdtDEEKbVT
cy6Jc/Pc7HscCUKJoO99u8kRSoWQKEeQIVPNOc22BWyACKWkiKq/yHto5C3ttddfnCPNAM5xNGQ9
qVgo5bgvQmTwRNGu3jsoEK9f80UVQi4HLZ9aypDrysp0X+09a9d6j7HBFhIOKzNN5hlBXc9stpjY
iEjN+1SVH8h+ZD6QREibN8hr79faNQVApLXCgKAkOcC5af2ygvaYYGqQMTo1Lmi/Dmbmp5kZJSbM
gqs6era/PtrIqbkmBS6b7ICxTvICOx95oyEId7yebczlLz7ERtLt1mu2wy+1APHG1BUgI+nxLag8
R/+piQF5MXNfqKkyoxy9kNg67ZQ3OtRWt7/SbBpvWYEC5/ducgo59A6Mq47PTkVIJzGqWi4rQU3n
uYavMEfsfvxx+vNokmRyTz47qTnNSVvMxDoNwbvkuGDrb61RXHAwj0+gTdn7kJ2vF/0OXuOyDuyM
0AW7aXp23QeUSSxBVftlC+v+gAbM4lUDZxdR7F/0f7uyC63Qw+sUbcBVaQaKi4Mp+bYW2ZEf1qi8
dF/TBWcctjmEddJMKZn699S1fFuTf6sId3RlSpV3jhNFE9aoqzKKJ1qKMSC3/dseNc4eNjurSPba
FxYj42ONJwD99feOY6fG91VIR6l6aZVVznzmOILrnd8m3JXL3raVJpiGM93B9LWJxtBVlnNJx0gW
8V+0rYlIvDi2RbPL0KuXh9NNfoMDQbazQ1wMrqH0LSDC5qtpmXuVH2eagI2niWVJdkxUNVL+w5Ff
+EecFynNky1kOUxA17B7mrI6bPMtqQE5LnCUuduXKkJFtxcd4YTxXvP2WBQdwyoeiDX9K2D3vMK0
Dwp80hZoG3BzxxXop9t+0C34LTRuKU108PKpSSBXXW5+IMra8XZU4lQCUDT3ZnOEqRObWd52TbJ5
NQkSN+VQ0Hg5/fNWbJZGugpbun643x7XTketfMWRzBL9bC6o8m8hyXVhJGRe6AvZmyuRs+yKPdAx
IUUPyxCjvwNVozMawkv+aPuzsyT+TGXKVxLNQ8sGlZDhuSHWr58Bz/yl3KThAWq/XgS+8Zr7wHs1
C1mTB74gwwK3zpKbzQAgp6pnkSoYjzUrXm4SUV++W6l46nmH6jA5S0QyYpJG/NP/jDD3Rb8l6SYS
9bDNJ0WDvJY9jz6U1yZQ9UlBWsarpVh37U9br/B8orwIqdzEGOso17r+4OF/eLTV1HlsMYJWsqYs
rzewz2Dndgkh8ISX9TqlIdzHULNonGNjGOujAxBJPxdKshhMkcXGokFpklOf3QVSsS/bkmt0BRYc
k+SL70VZF976UyvnsfxNIex53ckXzTDVrYLxmBmhSkleLnMYAh5HvOSJbwUUu/5Q5qbTPBf0frGy
TCUpyo/Oku51gBjC6eMIg/qiHtd70Pd77w5L0+R7ROE49dvMhouYTlHU0ROf48K7S2iMxpRCh2Hq
ID/5ctb6qereH+zBVQzhsYaeMPfs2whXoZTeIqH3IVQlixSROWCjxl3sylRRNrMdWmflRx4IA3Uv
t1pNBhy+jmFpsIEKTMRg5Yqjg//nfG0/OWI0dbucpBwP3F3+VxYRphobbM5KoscYVubbWwxEG8j0
nx1nQOJiSZuh/tAZn2uttBhHb/s42VER55HTmgXqdTViJIQApXD0FtoILgGayrYeh3qjXv5C8TfD
hsNPdoTJPOE4XxE+jmM7Zpqr+YHmVN9Q5zxSvwhngarZ3I9+mVE5E3+EsYMJ9d6hW+q9fakTggfe
SYihxMJcecJq0haQNCfr6Xwe2QugC9zFekXHmgP5NVdv7S5kfJDh885r8/WpXikVyjkflw47Sg5K
dvP1Py+yK6UulaVCrguKBBHEUKIAJhWhXsx1O6PqTlfUQoQY+/1UcU37DnVWJ8TXbRBing7WwZtE
eXdI0fYI9+RUzVMnriT0pLYUm+SorjepsDmYI5DGYVz1y24fM/FlatGf+X0TGvgXSE9dc6e7wsEO
wFYM7yBuO/1yU/XluCPUO/Et3PFzU4nlGpu6FtGIpbFe9Cr2ZvDCXk8qT62cKkVUJ2aWhane0lde
a8/B9YdI1r6hKo915rbZ9UYYYbEWklBFiTiuTzWch2v8Utey27d5KaSkfYfuwrStH8i+EdrOa/w8
sbzyqa6czkHTAyXhMm9F+0YW9KvsJsz2urNJeJw2eR9x0GVt4YEmxOkNHEQzsdtMBLv9Rl21Ofuy
hIa9jbuG8jLI4UMSUd7XTi7jRApS09N1JAo5pnFvME6PpyIMR66j0YK6391OpbLIrJCGcU68BFiP
kjbOUXReJX/js5RTY29JkRfKvO7FBmHoXplMRJ8DAW9ipSqyfGmQ8tQIHVL1mIuGHlEUPEc2qrNZ
zNeYdHwUDS7/CDsRGqXaXNT5fzgqRIKfrdU/N4Hw/vHpN5DMXjwQlR7Ib7abXlci1m9/nG8rRuBQ
r5l4Kal1JJ7bIKLFHdsh59DwntAaD9f6C9A9qXc3QHQzuf7Eo7enJmjz2ptZb8Cl7KepmpvtivkH
40qHlyXLovzkRjQF+LePtX2R8SCt2nuOPqrPj9SpmerKzks7an7abF4J1d8W9cN7M/wDeaJxKFL+
gNVV1xu1I1Uc/uMFyQl6UQ6b87fgue+ix2ZOG7HRqSO9y82kjwcvYOTZNd4FCWgiDwtuPK0JJSyt
h2W0CQQiS8q9/mHMCHG55Nv4suPCAXlhYxU9r4HeeLXyEym4FtPv90sE3LHJZ/PqcP+8vgj+ggTc
dnsc27N2qIt3IloezR670qdDkD3YK3B+vTFk0r5IWK6u5dIeEQB18CAH9ufN9coL7V/1AxztrqiR
VAxtKUd6qUjLGAU6mHI3eVsq19VOWow8ghboopyJufnXudxaJP8nKbfComflgOVoZokOShB9q+V8
C/qpVsT/C2zIFJRQ/rVvx5S563KXtvB4nS84XcKx/l/TAvO4PMoEmrKUMuzu4d94Lybau1AdkqD2
hduKnlM20u5SuZc7q9xQJ/l+udeaQ6ssZ9xJOtOAfnDDhPP1TyhVeQzVYTHRewIGaJ/7hecescT1
xsSQ8wR5zj4srwmx65I0QQVzp4uyEdDkm3JC+N7bP0shteXlBjwOZDj04oQbIcuhp5013hEKBaNN
qg5J97waGe/0BATq46nDfK24c5C3bJuQXc7FytLY7T3yInoKLjwiUR2tX2k36alMEwN4/kpQb642
V5v3saU3LxXi5trOWajkDRGhz9sLbqv1TeI0SPjcFyMI7i8OE3LTaiMMG3nOc9YDdOZ7CR/gFd0v
Bodw1MvC5D8XSw6fb91oj5jVJk80glPn7fHum3LtP8MyUufbkD95niMpdu+/XiDDMqDZYMIWrvcU
Go8yL5E97HV06zvriPVVYFEvmZoZ6uWQbTFc9G2yxu5ps9rs6Jt0NtlzANqTn9pedWmQt8rHuWUb
5k4Rt1MO/NTEK+HlTTcTcUeL2+PIsae2uE5BLhh1FJaXrYbvseQ5ur8VmAAedkqrZRweAI+s94nC
3zIysYy4CRtLjME/BihVuoGR7N2ARtEeO8EqUryAJS56Emd2uCoLAvnFo+xP4F6vatcv92wkM8x2
KVaXHeLU9r5itnUcXc24KlIjR99WDKJPpbVfqmmk7f+G0vJVvG5joJ30bfT1+cF/yEDHForv6MUb
Ay0dQKxYB/YXvBVS96lwaTq+a+M2cVu/WkqzNQ03Pee0+DkNTAxXx9vy16WwdqmPGRExRaVcQn1I
Ur9ayxfu6ZC91GVBZ8QnGrH24hioUtDDskTzwoYIWnrfLGYb7a8A8VCZ81ox2xHb0NyY0PckzvSJ
O/TkhaPck00rL5Js0k0PAk9kDmhFqo+lbpNvkhlu61ltmaeQjjVr0PwJ8iClBBV/NKCcgS/7u2ta
mnvBCnxJLEXxHbjp+6qptq1JlCjDbQdlK1NFDNbIQrXeTL/KDUsy2UrH3ECsX/dNY5j5GJ+HKrQC
vQA2XwvExycYJaK80xeeQVuDvFm29x3KpqHqO7FbtqHjSRTPQMHKcKqcy/aCZJnb8ObbgREA8dfq
L+wtzdljBUfaOdHwFRQGQcRBMG0gA1Y5wAMF1oZ0TH8tn8LtfWEVnn3+YIioBcrJJ8O+vV+VLEdk
jm/6usk3JHoimWu+BG3JXTKV9Nt6uyw5+9jxt2ZEl7KECw52ZPIDTuHusZ9tWcS5LU8CXI7TH1uy
iVsiDCTP/sMX0gFd0uYVmbf7jv5tYw/MJbphpWIJqWQANd0vO2iPDAQJ7TeKPd5IzkZhqAba2sMo
BQkyQ+kxQhOmVgCHOVSrA5h4ItHCFUPMLqeUSfOIu/EaJZympS4is+A2CNGsUy6n9UwUcToMSGBL
i2Cn+w5itrRJYuGDILgexHpBkQekFlltEp6IQrKfurcj4GN44CfYua4EkcEQnpqLs9h0tnU6w5Xb
gzcBu6U0f15uy1ZIpwx3WpgbAkvReynxQ8LRXB6dpRYsXFzkarycVny6lpcmRmINuAenPtxb28hk
BBoKuFsSopmJuZ4JFVV29d0OplZp3tUwlh193q4Zl+PeEGc6ARz4BF2gFkvYr/xbACleiyuEHbpP
7hOsUqFS1fcKrfBRC7ILIr/4y1Jg1lN4f8i/ctZH/jKwG+NzmAqYW75bfoutICwKin7ZPLgJrRre
8WHyAGL1pSF3m1yB3gmAle+tqPYw7hZqIPc40bMktkIR/E8IJNachtUVEn2B1QUL4XjEB5Y/x/UX
jlqbxEH4Tf0XmDxMe6HCX7nJooC1C1a65Gz5Qgt5Jl8M3JXDDOUuTb1Az3MhzKD+CbB+fL2h7NGQ
LgikInOudJyj3bn9jISk/JCkbCMlXsFItuYqO6REdnakB9rOomglkSWiizq/wz2LupFLjni1/thm
dP2kxHP0EmmCcQjlxo34LXM/W4fXuRBdyBwJdb6Ske0DofMVDZ+qdkvBCYlPWENy9Cct2/SZ8hu3
5GNtwSbcGzUwBuhq2ilY/Sfi9WIqnN8kPVPauuMUf5+WStQBKemZMerhFHAJ373jZiAgZuznvPUv
ODVdhrYNPjsolCfgNRZjH4JfJa0K8gYnzmGIs7Ci37EXL0sKM/PAZgF5AMBELcPZapAXSx4Pp23f
UCJxcKItvQ5lvsIUsqeymfNVagv7ZFrz6Z0ZRfSdi0/LSVdA6spa882XZ34Y/96diiCFG+KZf0cO
HflZTawH82Hua9Om0qYir4VPAa8VBtwPxuzGeS5Zwsn3w6YqWqLg8L9ZKH2rrM/hgsduJN2yN0uu
Qq225madS3TU4+sKyAUSdyMnhKX7uaYCcow7kHTxAR61ctnOzRtZEodF2y7lwk+PaM2ZJ2kovut8
7TSwqAH9fMHutvqxj9sBfxkgQI0l1IoKtL4S2hSvFq+1mtqA0XhINRJ8+nlWyw2pOdJqawXfVby0
nZONirS8iABtmIO9FFY0K2PPxzww/C0Ob5afClFQ98qTyfFH8V2m8p4AeL9zWa6UnETD/3CFqG/Y
uhHk9dv2+ISZHdqrbyrwvgOW8oxFhBCGejV1aLjFI+O/H/vK9ClgTpdteyGghQL4DWw5tUKKsvZK
3wBvA196wQFbyZWvdGwqRPqIOOQjqbUnPl+B2WKqHZs+V+yZcEK9W50KSnh8f3R2KPTeFvB2YpMe
0/QrjmkxzPtpL6rZe79levSIgl2AnTcKIjfMoLMXRMuFqvANv95337mRdRfKegqojAbkuK2DYWNY
Zdc+kvvlgSU8AQjlrn7T0LISxlB4RREpOhDclqYSo265f00Y4Zaijfpqzxtm2rL/eFDuXdAaXtxt
5t+oaXT9NnXClPwHtLqKsgt0RskzXyB2uvP0dBxLjHCKMexveTUBX8IxnCiwTR7i0pL5k7icDaur
M7CId96zSMStx5A7uYx9ksJUf6CgaCEPEUslYO+zjPe/XFc1RnaDObd1iCSv64VsYp0aMZKlMKPy
EgcDvJc8DLekY/CRbVUt5zVFp+SgKFn677CV9C8BgzC8TAHKgTBeXE6sySvTRUKbi3x2Ol8rSt0X
U5s+o2fo6rbRf73g5cBAqlj8tTTKRepSLfuqqLYFKOhKABmnKz14oa10JooZZucivQKWqwQDg2AC
xdJKi7/age3He3cyDZlDkXZyMZN9LrBtbYV96i3dq8ju4ZmEIe5tWvDTJKEVn7QzGyM6oL1huS2V
HNjSaKzvMDAgxV+B9UHXO5v+kT6e6C8FAWNCMbAewrG7j7Rxrds9nvdbRgJ3oUIjKXSxC22XS3j9
ETG7nuugc8SJ8dlcziN4WUhmQ2TmFN29ALKONMdMaqR379KnQEL0asN67wdzZKD9xX4MV+9ERbJk
W2ZYYVQ3mM1mrHirzXfRNd0IEYmUijdVEC/UVKMrVXccZcF0+q87zzZwUcKOP6BWSG8melmvXd+S
csUT5ifQePC8tl3WjXEQ9CtOzdjfdcT5AInZS1267ydDr4tZ3DoSVuzm2OraNsSen8enVla86S+D
BlnG0aFVvPqcPxgTNFjJsF+CLsV/BEiv+oxsjzNIv2BAAFeYl4Pdck6/YRdx9ib2fM6zSS0UQg/5
4HL5wSS2n9zBqikSsGT7EmGdFAcGJg15ooKA4yzNV61YSgHoQyF/FITbJCy188EuYq4Ue8/PXL8V
iO1wU6DC3WzbFWlPiWqk0/YvEJmwGcNTY5Rx7t5GC6zDgAW+NMFTg6rgRbguEP+RXzASE0xz1xBh
02HJspWIzouKXYsXIS620MFJ4CShxGlMFiqXQrBvJpZtUMQC3Dt/f1NyidwkI6COrxeMY9SUkhOE
mK8TMBbMU2mIw1c4vVdrwXqgeA4G6/PO3pSqfO88IYWmDYJxkwA+U981Joet8yzSWNsg1TJHnFyH
SHSowJtbMBZXmWQlvyltlg3erYCVEDCTymLUcx2PBwrN4rDg7acP9EN8s+XTs5kvLJyPAqdLAgtI
ED8lfvyxmNUw2NEpdgwLpLW5h6cKWKuexkfNAFJZzDuvr91kmONLSOqbwyjomq3a2te3tCa8i//x
cuLXh/Tbuzp3f9CQP2QD+gkMlwCbZpsuu4m/dmstwto2DAiwxiiceDgeCPF6i3ulN+KXivsp8kc8
oZmyNnprauCDoDk2yAB8AmUh4FvaD+jXOr3DgnHc51DzpELIX71nvUFlo9UXDXHKLlNb1cnoGSWf
nFEwqMGv9hrbb0vpa84BmNjsOcVRMcaePqVK5V6bHxOMI/fW448xm1iEmCy9bptdizd1LetD279l
IMx6p/9Vqp8bMsDdX1BsKHYbU+a0CkXnmpC1RukMpARPwLsKkiOidBI2FViBEoOw678imHPhyYKw
nFQKcSz8QCE/RjCNDJd5gfwp0ZBnppmJSmwp4cAMwFnkw4SVIm/1AvIu7jqOPZ1dX0isJDFVzzuy
W5TbvN2NqKbLtH7XC/6hoE91QMWv/I0rITR13J9zdmNvl7qcURZMnkKfyHorXeWeyzZUJ3MzJftY
tQEvKttF47tKhR+1SburBL873ENdtaAd89b+4rt6iIuTGx64u1Wfu1RN2XQ+7cTVbMnzIpyFUKxm
rXU0LFNvXjl7F+tbV/O4B+npQJ1jIcKe5Rjkb253u5+YlGoViSPXo/rpBHCqLnuSqph9pmTZuhrA
cxBrN0oF0IskKS3pOZQuMw07f+vk1P7zkxfmq4nk9XVKJQI6wrTa0Rler29Wp/n5KHybb3XknXtn
gQ28mqA2RUKl2dg+saBMOXG0XbiOwIHm1j1X5JyR7ORrnuwU4zLQrHkd1jexJtrYQk2CSW+Mw+cR
zYZT9SdEhrzbdsiyuI+K3P/0jtSgLV6PS+/Sywi+G2hamNEIfOVO8v5q5HeWuu9/SujHTfg61BWh
0mOidWWTfldEv+vvPCFVIqc8FyJ/ZNYrX6+fAv4JaMXXnxLyMcW61Pq1HF0xMUCLUqOZyesMW19X
uZK3PJg+vm02ihlg/0tTgphtlx7lQ+yTLMdxm24skLZjVHrms3xRoIAo6i7bRmjMN3UiA4K0tjDD
CzrWLO4XHHcNy9U4DngF7G2UnJdxTqglGV3WSpO7UlgsGWrrVCCTc7W6pOfXvlpqF4/a5FZ4+Y7C
zMNtU9CKGZ8WYP3krjQIpCTaaBEV8PXH+TNRAZ5h/Ppr+CAUTYl6SV5aXLFi9qPg6ZGvZY0Fxm6R
y5oAcVlhEOXw49Nw4sMjklm0bay4MMm96t4stblbyU+ejwnXCNEgg4hGRsQGMR4RBduhjr8mWl9W
2rVZEGbYip83yDEAnBPHKCAhpD92AFqMDtzqfFL8hgVmBdaR6d6w8LYqqbyYI0QMasvQgvzUTUmi
eY0nPpz/1mj9+5oyMo092qKwVCBLMXfIp/ef7cX45UHBOrsSPyOmpH+rs12u8kDj6yyzr3f7jSaP
gNWq+zhmSJQjuAUXWV2gcCJDFlCD4yrPoNWqU6cLa15kZrWfRefdYsjp3a4hXgSTywXW70jngZ/1
rsZ/8n7BzP7Sao6B8lzit1Rws/3NaYsEsMkHQotCvNuBRZDDvvv0AsvN0ZkjA7XmVrxyWO8pRTs0
Q+UKA/vPqgFgHQw03QcSY1/m1MwVlj9f3eSs4Y5U0mVwC2x29lAzrrygzpUA2eKc2ZjCvBK3BXCF
x8X91vk2qu7V5bTwK+47Q9GCVHi+gEO4IZWPSBMnFrj6rgkUxYmiDZs7w3Ora4d05YiN6SgUMCWL
SXxSkFuxmDlOhPL4r2G0japVkjF6dlapDMfdkpQhMAGBrinrM2qCUU0/K7gooKd1u1BNNZSjV1wS
6YLmVG4DSDsZc1e7x6WErWAH3up4OXZDgvy2Ey8lENkagQ7auwBSVp3JNtkYRA8AAOnoTE/3LGIV
lS/3NxAJnem2/jRYNnUNDjAy9Qleil6dSOuFPLubHkBriv9EWzIFv0pvLvGjo/CWWLUgfLQidemm
UTKAJqcUuVSBmTRC6yLZqgmJYKxE6IuRw76lUw2kaI7ipkq7nlS9c69YlgEXpwVNta7QqJCAdU2l
vV0CncUAPfNnT5fMYFQ2OCCrGYpnXzA+IEOyJ4/KrXZvhS1wOVyxAqidFwucgRE70ndjf0YWm35s
YdEfZb6p/gi/qEkr9KJ9dHVEAQfGRzuOnSSpJl0ScDIyL7HFkI/EW7q8lupFDxNU2fRamF09REPJ
alJH+IqKOf7pbAlvRpCxBGziVg73e3yw3nS38YSJqaa2f4myD9uFtVj5sMlcb3Gv2plcdNACDndH
LbTj7mtOuFiFfl3yAqN5qS9Y2uSyuyxS6qY0wYNzq0Bfy4XM49LxWjFuMimt4uuOhv8zMSlWicza
wBmEj1Z3Ch9Y5GbO/dCqktVcvOcaxA2GrJDRz2U0rXYIO4wDiV2IFRL1FBedFrIkswQZpKMFF9oa
BKZHTdCGh8QaCSOvMeaBqjci4oYCRkT+/KrYYEJFHisVjEiY2ztDjrOiONclbH5nSicanUkkpM6v
zizCwhMoZ7x3Ou6DjtYQDx8ujk9wSnh+B5Xv7q9LxbiKCv0lbSjgGIZhUCLkOgZWVFQaSvtbw18e
f3fmT6TGk+9MWKMl588zNB0+er/65Ngq3/zLgraSejpZqAK5CP9qX5uwP/VP/GMuWYG1bppfoNyG
XWAuZ/BG5BckDq4tOft/NesXChsVOVewEDWcpYNmBbAVmY3+NYTnyqV3xi5HuZf6M3pwpYWKMEL9
3yUP68NBeKWkLhR5K0vURpbgVLKdR39SfI9oOnAuAywaeevW/IaFRPAlYvovxVCuJ2i38GLuhTLM
KFDS1ksLfQ6Omvo4RhRSAHDK0Z8BJovPYFx14qawT7bKlVsGoxra/UvNwimNyVWCibbhmuhwJNmz
8AonqCnB75D5Nm7AOz2ZqsbK2FracerVvvjkC1OR8VGFffoeT7sdV6uheCZoYAg0UoChdBmI6mke
0JNzSc8k4JOM0gyQWQJmp8O8BEslqwTsx2pIH+hPMNB1HuybAfohm/AVz3zt5LEp1sM3mZtNs0ey
y0siyK+4o/MEQZolM6F5Ols6LUdFzkDZAXpOSb3ew/QhrBPwWHxbk/HDuQoh2pZI4LGzkoeoJ75k
0psrCGA0Dh7GkoIKNWy4hHs/Natnm4/w/0WkOap5mP98bmS5Rbftr2NQu1lduPj9hRUQg4GHdrKK
S8IYNOo5IfXdBQPRwyxthLNJNK+9Qd3GjYg2rcTZWFtBnGp/I5SdDYci1td+R7a4Q24dVv8LGdoV
R/KlNJsxcpeHuJLfdp4GZX9BeSDgCnjdYXUFYxXwyaC089ElbGijDoC3cLAzhOFxPhz40wKFgPBs
vumNrVuwGvX7zGtWO9pWs9ZAbEFykjAJ5YZDFBVqFp0YsvOo0ByqF8cjSz1Zq+oiykDWfW03jNYi
FBU4U2Xxo1wKcbZ2/OXk6qRtOstkUAg9XdON8kAstNkEeKr1ABBjo/MEjcJR7gBhBj3oxF5jS9Fs
r7UIAVBCdwRa4ytWI9XYKBZ6AUNXFNr2Q9FlogD1i+xeYv9a6HlmHHxjFYecP69HmwPTsAetKb30
AMKQZVEAf+iY+pR4L/ohxDI9utqvt7MR52NkpBBB3fFF+K/sOt8i26Dl6TTOi8EiTUKcZ4ZDzmp+
IkXgmLNKxcD08n83ehxqJYsImhTLwZYVF8OwBmldb18XgSA8D5ZDhPgOGpoCD0w0dEMAzVRxUi/c
quus+x9crgRU23JOTUd5zyqj/uHqtKYkQs1PoEoY+6xhZrkg26YdIToualJYtKM6onEb3ynZyhtw
THZ0Ie1TZplUYiDaGakD/aSg0oxvKmqeWwsCuhBxGqYTf1ipLAbZoKXNMwLghMEtSAl9QM4pM/jD
Ew6PBelhLrRblXexpeBjrwmxfV6W4oySk9yY5Vv4wS2n4DiJsMYWeqBys47RMYZ9Cc8WdA63jhnh
a9wUXnjW728ADaSOcHe4oGH/Mnl2xF8jfeVBmQDk6xcmrU6QPQiYpOUkWOW1Q1sEkae2pVFO6cCQ
ovBTWRPJC28tMeze4v1WfwhbDd1K5fk4LdkN43KTLvzkSNHLzKQS/oak2aZREyxuK92DE8Yt7fxy
vvNMYKzP79plcZdd30QlD4OYRdq/B+JJyymffYzAXIcjW+wWsdgpf69ANJJ1Zj2pfb0znU4QuyUm
9V7HvHEchyHGlvtJjwNH9C2F/JY24Qqq5CP6VKXgC2uvM9S8tE2fix8CK1V29kAvoNSG62BWGNSq
zomfb26Dc9+mnRKpawaOEHB5S/+ouFtF8HE/jssQqLdDJJAtgAf0u0AcwcQJA5IEj7VRu2O/jHJU
hFYoluZqaPjLvpJmRNnSBEpalO3VM4qEfskBaCop6VMVscUrrfz4IZKy/PNl5dSRdADD1g2gDiaK
M6Tgq5Y56l+DekP8JwnbUP6LIH8zi9jX3LFoVWFfettiLuPaEJ4dVTVkMhnCshwCXysLxrTqwzSH
+vjkU88NteUs3ONg4o76v/a7ofKybOGRmXflTM0T+jk0y/5enMGJgHZr/GbbSlKvNIoo3IP+Wwvh
8fpyjGx7tl16QxGTGOlbE1A8nSFSHHrv2Z/ZfMKn1qpmCZ0P6ro9Nx8C+F+2+4UdUHAYwRz0fl/j
FLc/GfEMe7773I/83MxCMg6abR7foa3o9NYvfYSd5vo4OjysplbXPsyoV2jfwxRFlY/pZReOuWzM
yGiQsiZRAf76AX9sKKPWZWaOMfgZ0t1IgcIPIkBN3Tvx5WlaCsm0CA162TPPqNJkVoM5o9TpdH13
ZumAcnkeYppnEfOGpr58KacX+E3ElgpwA4stW/TDUPb8yjAFBMq2rl5CYm4IplMie/QTFOUhKJHx
pcv0xz469H3ZfoYGSpyqDclGCgEe25gR5wX6Aq6C1E9GpqG8lL8ImMLB4v5h1SBY1hDTZHLV4KnX
g9nfm/IEk+bkdzQJ3n4rYu1Y6h+J0TC08ppqC2joojkSvYZguOZBfho+lI8nbz2Txyo8OKUjyedV
MGVeOAS5GG5bJGWqlqNKcZ0ZnNWdyT9opUa7wAxqVGRs4/xDwJ6ioJbR4SaMXfXzIJ6njdTbrl8b
tOjhro3PGh3MJDX4zlyFDBpYigNSXuo5NfzqkDdv5oNPb+ATm4imGnVpdQHqB8+FcIURLEQm/khg
X+MCIP7NfGSwqdvBp0R2LcMayknL5K7mIf+uEVVXagGlOKKOMg9iBK92rkz3L+adraEYRrUyjWpF
kDC1bPwWFXw3TNAkeoGKjzxELM3sWhrv8W6n1hkw0UfRLkc22SITaRm8143Aid5SVG0G3TznJK/V
K+SV+bdZjqR6LzPJZAMjx+QRXl3FpEaWQpk0gvogm2+TtBdSO+e9aGQQxXD852tYZurI+mF3gAkO
ricFP3bSs1YomYqapgWpk5BW/H+rBzeJKIHOB8xWRDW1K0cWO1jku9+m5sLB0H8Hc/DcKsXmbss+
a4eDA7Js19yZb1y27AwwkgP4U/fxqn+P4miAty+gCiK8QL0UIHfOmWYIMlABV3EFa70FMO4dggRD
HX4ZEcLMDCaAIex5KftCxY/0E++yhJCTrEoCpYGX3zT8Zxmt+k9Usv7YbaVdKHocAof9Fnkvj3V6
IddfmkxogwZuCLp29DvZUftBoU4s5m1CXvuHdBjVu/xjgnkPvTchbKP90AjSdM5XvdP/1DRdf+uQ
JbaIrrbh3Spo1rJ11iCP/+gfrnp2qAgt/WgEekpDXcB9GjwX7xX4so1ww4eUQ8Nw3qPIXJmY2dY7
GiNGd1zHa3/yoZxO6jHy1EEVyEDM8ibqDQxeIAG6/alnJZQy7HxosRTY0XX5YFGCX4a/IaK0DKDz
SYJtVmYKs4YgfQXix70uR8w30FAfZaeEGoADp5j/m8lytQLsxWq1y5hyv7knwu1D2OO8EMr4JSFa
Wt/vKJwibkE+BTdHVH0zT44vQyY12TOEN8fxYsgng//oo+LLVOb9F9N15sWgAJ7IMsR2f1vqzhAW
fkG2PLTqAVoV6QjfB2O2VAczg25QRXE/BT42ZniGMklCx0ltAgTUS4ubOxPpYXVdP3vpHvsN5SfG
Vcsn/UQBAJmpxo0Ygpk6tV/MkxObRoOnSD/JP/1AXuWkTbkytcDu/VBaaznVBiIPv2Il95+dSUPt
EbdY0uKiERX5kQDgSC/kUpAR9YzcyLw91wbbRO85N1FdFDTduR/8rs1DiaHss6ygp8AW2RHmGgo+
z+JZ/59oGoFtOpwlYzdIw9ABXt/GIRYyQlUs5TYpVOwTcqKNg3rP12mJYSvAYJsLcelaYs9tK5dd
bwLqdqktjLitNAjw5fcErjFAzEjImlu6VJIjyIi9XCVt7t5SJIxCCkWeWqLwkPBPW2vyPu8SM9+K
TF9SvsA7NorxR/UBOv/LsGoKEzuvzu7TNM8eqJ/OP/nMcpDY6/RIuGeVZBAFb43sf2uJcXQllaTO
aSSymwKWoudh9Qq4Y8AUewC9RfwDHW4z7vjGudjgDra7NwRSnlB9MBKSmxu1bL1yh0cnv5KXW+G3
xnsY+TGZEr+5nzgyTeTqNkxP3UUFQH4EqJZhzADrhnG+Iq+d0G8D0d6+H6OxoceXt5iFU1uI04Zp
qS5Z8BP/cWfN1b4hBMb3X7dhrB/zVpzc0KjPdOvWbOkS+g3i3r51XvKOOGYW4e2MgIy3YmO/tzUs
CVZmQeWor4NPGpdIV+njK+lEEwnyRgoeeqtczaw5m6IGEP+rjF6jm+qGxHdslnTCQYG0rC6AwkgQ
rMbrMIWWCGO6T6CUc79G5Nms5zbyHRtpbpEyEpE4QweTa16yYkL402PyH98KEAatbAF/XQuHmt38
5Rownp89DaFR6FCC+32jdwKCvovq0UJKdiz8L1uQ5aI3zAbNbLqbSryZPfBqtrdb8+OD6SchtM1e
vbBvlkEtdAR8zIblycoZdxydh3OE41zqTRKm03q6bgs0G9zD6Q/GLwnzOysm/a/GgfAexwWfWBuY
lCmDfDRSoNshjWEl+/fElhW7rBQs1Tza1fPHtL9vGV6eTEsxlpkBTn7n6HTVAjFKs8fphoKf95jC
kdqPZbOQOvdtVO0SIWo214rKfTH+JNpB+zXKOxxAPUX6b/E884WB46nBVRwkCCO83Kqmep3/I7XC
VsNhqwA7zvJ8+qKELGtxOsJpr0vXMNHKjDnp/UTyzpVwu3QGqNylYr5nrd34BNtdKSP0gDQ9n27r
CKsEQnGrDf3yzYz8txZF9kz2ksKrt1uC/mP/r1o8m1gdcSrmBDCLcKVdODqpC2Ruo+US7LmUSCBX
zMiVpmxh4dEozqs/OsYJEpiqOAZkpNHXNHSl4pagekthsA+TxOGiEWZJ71QVNNI2VeM8QTbmllLi
yWx7KXlAvF65pxGaIgOJ0c9P3vX11BihvYHlrk+Kjj9PtqcVoCxz6rPMMpXwKBFvKwF27Z1O3/vN
m1/2DPk6YQqof6hTyR0iM+NIv2B+d19Wp7HueClGzMcj6QL0C+rVpviNzZQND9Lw/QcNXhMPCHV3
DPUw3LwxvbIyrOJEfln2qSn30t3erKhsWVnPOvwx3FQOejHpmlXMKLSIXZv7YWSfEdkv2LosdRXY
8llEhzfFkJPHh1z+Uxamov1VLy9B/u49UTa6rPBhkcxfJKb5gxZf0UVUmrU6C43e7XXGCzn75ubx
o8e4Pwl3/VYxJ+PK7jOPzs0tYVxc7BLhhJxO5b4MO8AhdasfKFt02jOpLdigU/szhiHoIc8v13db
Hvkb46uVkgBu3p7cY6LsS+EZsHbW141iFchOX30zhhPkREukw2xDkJbL0LJZ7iKeeprovK3BitqF
a62FBRvBZJDRvmvKv1G5L1+iDQfVxtBGVWmRsH/lKaFKGP58GmnkD+ig64GIDYZLlLoI6B3OCoNg
kgHPy6pZznIXNKSoHYJKSsi6csVM/1iTyYjNEarb7xySpJSqHKZyt6EHzYAG19DqdBQBY6p0JODN
EgMODc+9zqRmirjDy84PNpGHVqSVyQSL9yAnrQ5EZbvXbgA+b50kVONxU3gEkyEuzLroFWdU+Atx
8HbXY09z22z+wwY03JXZzjjNCEN88WpbVySveaH5BPCKVG8+BfSQcC8AUcznVZaLKubYhfFWp8by
3Upj7MO0OD5qfaVMkZaJ+A+UJhYrIKL3C0npQYrj3McoaGc2bvKgUSwrFn8iSkU60bDgrahdO7xK
wmBl1jVzQp5c+RRg6avfz9gYosJjRSmuX/AjGUSZdcfi6CbcggzIEe8bEwzL7ObO6zxfgkVrz9yC
7PofDfKS/zr93WgkSKSrVHXyp2RwCRk8yU8EI4fYPMS5sSiXjpIYX3cAnYiMnaI9iJ+cSXix6Rax
/s290EGGD4j0PnIoOZLSpmTFLqFJZaHUl1LtEg5YRiVfKvGaBMm20cgy0y5h23rxcFInaF2Ar80q
QdgWM2Qa0tIZkQgxuiCwZZPqj/KTXyESYq66prv7vjdsc4ZtU+MV99X3QbCWnOk6b256EcaYD7m/
93fjM2aBw7W3Vqsx+AFOmWDjGqEaXLABDFjYSoDpVqlhKTu1F+XMd4Ov/InTCL0LNrQj8BR7w2XM
FooJtceK4jF24ONGfY9kYkhlJ8W9njJ/Pd0d2Djdtl64NpD0y2H0c9gh4n/eQ7Y27GQ0Re4U9e5j
ztbIHI9A4iHlLGXFo/WOcAi1UTLdiqJcNpLnJbRsC2Mco64dwZXViCFJWNyaJ/WsQsSEsD9RstRP
+a9pMoZKVoRwQTQYM3hssjYbBNW98/65tycRz3VGu+fobSWtOO0GoltyRp7NX1SSWiljMndwZl/q
jrcGAARVnBDkoGUZ7lZTGn4ujrCNGCbjwp7jw8P7K0HlnIUAey9i/mXtRWWuFDnY4yrSmuq5qczV
Xqdkp+psvtXd/PD+juLWauRVnRyrb87FLDjw6x57BDaMPf5UZN5LLntSiozNDfLq8nH6kdcETYyv
SDpCLHM2wD7gS9Vz4wbCiH2CG5iVY8T5okCiHQ/qiTM+3pz8OPhog63VUSymm1iRHnhyuQbGCrL1
hea2TilcCGqSDUcKt9DU2WUu5hD+byqcdhl8PT78nUktMwYDR+l9JuDjYz8LYGmAR/OrmOrYEjK4
ow8BZLFt9LdHvzjKce7HLXUVbn9hg+4ydR2lBf1DrGgJlO1Qxi39yI56lcU7lHzG3116uTJOl39z
LsWvCyy894eybEy1qJaz9WR/0JplY3Y+Wcm31Yy/hbXgiPJ0WaVpJYI6edkfDeRwWVDoSIDS5Faq
Rr50Uwh8XApLPb/z8pGhiBehprPCKjRLCLbxzGjwLMhYXhQc0Na6t7vhQyY9wccWhiRoHly02Gim
+nb5dTpgN3NpOgsSv9kH2wD9+B2ul/4efBBOcW/bWtGFaEr0Ek7oglS0H97ad5u3GuO5LkYWnWNn
R2jKp8GbyUXB5GTGQlCd0OL5qUu1R2n65RRkITU8egIXahS74TarMUPLfw1gKAZITGD7np/i/bif
geZdEF6yiEl3cGUQ4JRkwRxODtWUTkozi9qzOgk5LnX2jTLnQzpedshrgn79A7L2w8Vk/38zTk4Q
+/2XklAeXgAEqBPXHsR8uZv4rBxG7GKU1ikf2FJAJt60hFT3/w8Y+qo6sT7DEbUzLK29SolATlru
cIuc6XyN0iua1T9+G/WFLQtIN1A0Oj+fl8IEnZ4q9d/iX7yMKdBDW3R6CgqISBym8eh0R8qhdQQ2
mJ0wT6cDOhSsKlCRmrhXuJRUXtuVA77b5W/flfJxNCb7suzNZQvh2BFYse7WQnxSzr141u3kXP+T
HXhc8M//FiHBc82QYf3MXAlJz6Rm247KyanZ/jlE5uNJdJfYnSZaIokdb4RI+Z5a53jGLFkWV+sk
1c/Z39KaZIlnqCcCU0g/ra+z6lX2czsbuOe9OklK2jqGL/+ye1kyVFMfKtKDhfvRg+snBUsVlXxC
8CzlncQHgoBq7P/Y8nciBW04wKlLc/s1caZavtJUT/OyAp+7YqCT5XPaaJ2KldnZdgik1+7mQniy
qXq45umZ5t84D7N1obaNZNAg1cqerQUy464QUmx6Kn5/3cLIIxurRsOjxaq5SyYHxQ3SgFNciF30
B2bkES3vsbfvZJuGetAwts6BqN+CMlP2x453wgEOSAMj9oHsJ7fAPxQcAdOj9SqwrF7GAnExyCHO
+bngpxREeq08N0h/5UtbTW9G3nzqGg5vh6RyNrwR1U+fd4vCv/qi8EC4P69M6mO4EmgY6N4VzWBa
Y8uS5ouuARsdRIDkG+iCkyMW0sZOqtIvIYtKrOiH+/M6gvKToP2gQJ21SqDLMOUHtgAwc+hOdFNV
pSP+Xe/R8u+MWjta/zIRrALj43GJpfwM3ctBqB4yc1X9a7uRwMe/NMYx4fAfbOrj+LM2VvVHwcFn
v/7sPdmAX/fYkCF0txfiAN9hOGfp+FUIVq+rayN/aHXXg+NBHjA11sC2+unENzM4u5x8ua2s0sUa
rvUmKlyrgPyrIxyWjRCCSFXVWcBbQRG6VXvsumSI0f4I/N6Ygu6pL3G+tTtQ0JoVVQ7EQZoywyP4
fZM0wSoki4k66Lw8R6DGJecc3e3CUKHeX8UnFcy9l5Is8YNC31b8pMRPgOu7TglMIemhzHtKo3gr
aQ71/xD2BtIP5yk+7INNxC/GXQCDYKBqau00AXnjNXgGb4TLZtrByNfHB2KegnEZxc4tCD19/udH
rgxrjnikgDm+CFFEdyCrlhZ0Lqz/9MPBSosDa+kNL7C9ZN0Xa+Opl7oJw14tM4zbaAcnhgKWoxhk
88m2/XoAS5yaRJ/HagQHZ+EyFS8mef+wGuM1XH/BtEupC6IDQV6gs7TI1NvvdhCnDkl5ikAQYjZP
C4DnrNBDYVo7ZjmMtvuIl94/TlxvH+JUpE+UE+wzDKymgRZVDQquCB/2OOpdTVqz4BamxRWkjkSi
v0B72/D/0/gw9HnEo7FGiCoMGB/Y8RszmaFx/JLY09lEsJxYevALdNND87hlB9xH1WDd6utNZFcD
d5GrTJvW+giuh2Ve22XQUj77Y7Oc8l03MjglCBjvzxPnmF7OYYpN0ytpog8wk4icVtu836y8fd+5
HnN5bBakDrY83CBahBl5pfBVcq6egUWZBnzMe5hLXxUkZ0PWRV4v/vibQ9feBEcDN4iY9oGiZAiJ
Ai766SSMncWA2TQFQYidyFrqSEnoIbAPtfoYiGfkNoDYsc7TESaMTloIPP2BR48kt9HWoYJ5+ak0
xiqbYTlCDzD43MObeCZFO0gHtvC5kZC50TsjFOBVolF827BgHhVkRA6VRi1059rNAdxqfBnVeIyF
Cj6TJUfe9UdpDW7psjLPzJzUSHONGD44PMcGJvofz7GlXF83s3UIlsYH9vkR18zy5tyE9a70kMsR
i9ASCvKCjHbTU/O42Vx5a1ZAa5pBoP54vq6IudzhKwfN/CdewHj3dghryZ2xuW/x0zMnVXzo/BZ9
Eqcs89EzgP4ZmT+5hAJEDMyKoy9/4yXY77r83KFfHnOiZTRBM6qZzmlVGH8+J03CEu46Y9aMD9sn
8e3HrqfxGHLZuDAhHeamtYIbM5MoMNESALyUQLSNfF9142uFG7DbZKbqjxRYQpzLQwfydUqJROlO
ERON5msX7HojvAFhmSJ4Ug2fwUMoAvb+dPKjGDf83xI+C5Tc61kj5YFYWZ/w6ZFuxgRk2dwJRRv0
uEkqCs6ySWtx7lSFNjqgRl+VA5DdRwqqIcJr+YFI7nxPSQEmUQmZBeaHUnjZpjpbnV6KxyW/jveH
UH+yW1RhdB8vmLBmVkMEiosfTmuk+D94CnYO5yXqqV/iEx98vKT10ATfDO198Bk1dh2fUNp+K+VY
M6KfO3jPSQyVizphrg3hNWGtUU5ylNB1cVGvkZ3526eN3VPqymj3iM78HoG7zocFMdupB3uwFKLD
rNyC1iuevnzY8Yh4J4u3r8eK0I4NGt7DwdzYvpyhwEB71VM4Vpks3n0Z9YEqzRK2wiZUHLyLQJrs
lU3+lL2+5aIn9ZQuXUocBgYHHSOrbp0dyHNoiKLl6xghkeTAFmhd1FdqZtU0ori6ZnFilJwDey4a
Y5hwkyLSCf0ah+d8f9GV6FTbnHWqoT9yeAgFRnEuF1TVzkw+YLueDfiIu1QmGlZ9IEzc9HqtEbD8
Bp/zy2ojrbWvEgh2ng9EDzjQktVlABrVOQO/E05gf0HnMaVaVhhKk5x7KdFzQFrAp+vo8u//tnPA
PaYlNMo+Jttogy7+FVhqzaLfSoyT9ZW4B91QZwxiiYJKZb4H1MoJmi4roM+qLQoN40g6jpqjgsPd
eKHB/H8Tq7oshVtHu3dx4dFxI0xqjTGmvT1TnvotpMiwP/Od/FLi5CUi6WFWHs4uGosczbuIfXNP
yuS4U41OBb8aOZPzsW9PjOtoBR/2LYpdyBFXpodC3afGlccRyUmZTWWMsLVRXXS9mztMtI8RGuOE
65vL6AmYaEsvqMWxTgRKN8b3t0hWN55PJTTAMSP/8Rn2Guezasbk0t3VrBoVVBAZhxGysvmY4n95
1A3TNeKXRd+/l70moeIyZdj4zm7XJiD+XtZZQ9rt3BT3CJeUQVY+ub7HoPkbGEIH/1BU7ZnK3Cgs
FJS7r4rkJnHk65GcqprqDCZvHUWy7U7dRQrRDiykArWgLKts/EEShsIm+dEFVpwuutuOdMeCvXXQ
XmmI60PhoBQwTYAsU/0k07CxRZS8GXElVgkzp3ZVBraFoBhIT7slKfcdcFjtC88hWSxGGVC1mKq6
c29PVfiglA5uGQLepYmOoAdSXx2JEPWbOc+c0MSWsMIz8PsEwIzmCLmj3bCte44XvXRJv6CDNbtq
AGKmQ0hlVRr4uBgzQHK+1Ry3Kwi7DPlyV4qHAudmAy4zPeJjexCBRilywoxAkOEIhwsAz+nUPNqo
MiN3xnf0DKchCSDXYR9nVbf+3nsfeZU8i63Q+ExlgTZuIx58xDeRVkvgmoT69x6PzI0b/EwsFCfJ
5ebmKIcatsan/qxT/YgWg9Ck0OAeJuwpZ8KcQTAc4wAP6fre0CNCYDsFYXUQYzNOrVHQTbyTIh4p
UkskuDf4u32W9hs+rKRFJqTfIpQumSTTobakqOJ57ALvaGTEVXk4Z2VOM4LKFNlrRzKTpRx2qDIc
FTTkC2kp4GZwrCpeYYSCFieHtS/dgg0HPBvC/OaK63J/QG9zqS4t3LnxcQ8CXIQwzRQTjZD4S+tS
qHD47mElY0/0sZq5HFB1C63cwUCwBz0KPlyCDUJXLC0uJWd+yuqT1PINbuB388mF1WY7R+hOQaz3
SDe3wnyE/hfW8vTqE/lHSbZun4ljgRBnuWXF1kkqHFhRDuCV9NNv5mXaiK5TtCbDyLSO64WtwPPF
WAXi8nnaEi+hAWl72zyZwLlFzTBn+qwpNn5+z/00+EEvHhDyK+d5gcTBjUefJFBFIEg1q/MlU5Ev
8RXksoQqgpNpUVFboOjnRbU/fJBpbpG++UTOBnAk6E+VsAEAMnXcDy0F+0FqGgXhxgtNn1ZEfRsC
7Bj2vRc1Iw2dCaU7TXOX1aWQeZqWtFKAH9nUkWn9cejkpRVlK/2XpMpjig3ddj8jxFbTH90x8HW2
f0qClpHT4lV8jcDs4/nGQ3f6gSVi3UfTnHK/YhOw8OLlhWhp/9lrowSGJzHPR6vLSrqA7bbc77kx
6lJuUZFDfiiLJaM72byatkw1m5EWZabLHCa6mINaINO9NlUsMIZ5Ih61EOPSLyTUbm8Y5WpHBeNL
hrKrGVbILNoA2voGti6H6Ipst5F4piFD8VXEkMDz6YrqK1jKVDlkusCf7eXhcyug1GBl9GmOVN1x
rjjWw9BWQuTlBYssuCG45KrsJE2sad9f3j+88Vu+d/6d5nFXkRk6G0zXCovYKVG0OzRv/+6m+Ei4
W2NWoai4ff4A6zSNvjjiqjvqQiRXk/Pmn/8oULQSZ22qCe/Q3LQL5KWbZD6v4TN4cg+qcYASXcX9
m198U4nQ2N7u6dX0ZmbVGCFW/aChuTkkt6N1xnUF6W5ZpFhzZGEBg2dfygbJLJuy8oWgMr0ysrqx
92UsXXA5zgtU4maaqEFmshcgEBx/tfObwCkg2QWlZWkEuaKIq44elAbP4yz+XyvfCWIajTDi9KUm
+9UZZ/BGHoDUIsd/m5eR8/itLsfPss5310A2clZ8UxFgd9yYbh9qz0ivZ+fF6gFUuf7gJHg1nueo
isoyU1kknSuoCKSI57W3xfOI8bVsYXXA/wMdSmMRDwPxo19RWhXu8wEgH4KJVswN/PfjTxWKc0Kf
C+buIuO/2eYzE0F5qQn6XAlj+/G1rk71KZvkjyq5hirLxxAHj18PLw1MDXllBI5xy/4LzxYE7fTl
yrIj8ad/N4XtzVNd1xrqpAASrDmkxQwdjHR/xgtFuO0eJVWo2pK23XeHd2c0Luwr9+mX2UeJmCjE
nGl4nvuib7l+aeGX/MKbu4hboIwTBY/oQjntrMkic8JfwVlidEVANekFS3+v6Yl4troZOjCRs2qj
ZncQ8yPLPoN/RiT08sq8QUOO/Hp03i0xG2fKWXnie8b/FaRE4mA3k9T7XbXlzGMphlUkF0KlLjLB
ukcMyDtR4HbXyu6kwwM8vx7LEKBQK8eH3FszslIbmGDe5KMOgBAcV2SbBsAwkMJBQeZugDNBNA8o
0Aym9YAMzXJCwmcvk4VkYygf+4OkgSiQo6DKIlV+wW3NFKaYS+KmyK//KraGA2W3249hEpkFqdJ5
VCs2Vmd2ZX0qXIvxqg920vOwdq7WvqAbu7aDauPkc98G6uQ+VJRggumLJlxuaxF8YMlPGF2yHarp
1hL1DQcjOtavrpiNm2M6skxMC9zpp+r2z+OIt92g+BBaLUr5FeVVApLmjqQT9DXUUVRtcdf7vzfS
RjpQZ+3wvKfh8NZzJbTSfxNzzs1YNiF0167qQ73cDQSe/qix1AmR6hDqvBfvU+yFOw8yJKwRRKTZ
+4ojr8HMY8nJFX+MYh1W51p3Nur/rVZFLzlYWSxc7WshN8tIzMk7wOOsfVe5dV5mHCgqySOJGCjF
Ad00jOrJZ7t1HubinalUoglh7JWOsDhMh6uFOsdzqaoFk6F6RTQOec+UKBB5UGmJMp7v0PhQ43eM
D9DRih5+ghi2RkhZhwAwCBvGzseLJ7lO73LHyavubBkAlHhncoeDYQExLp6TIqPHg+RISCPVRnpx
5fQDAr+Mg6+shPrsAkiLgTdun4aRK0gqnDkzqk/8u/Tce9DRu3ruuU+HeCaFYSvps4liM5zD0LLw
hx0Y+w2rjmuAw5jQmQaToX5SKecO0Gj8HTPi3gE7+052NGm+TzZ1BcdrdKvXrOwBNiwBjH0gcoOz
+dSz8uGiRqOjPR45fVttdsHqTK25iCCcwuLFIxkyQZ/v2vVmUPYyAj+OQ1+9dCVWrL2UD1DwTqXS
GiRq7o5b0eXQulD6WAzLKsIVXBg/rMpFtmeJ8Z3quE0D7JMN5vIXnEFQdhcJkamgAzRCgUuA1P7k
xyyrIkxlkcnRae/GRtWJ+dmeDixE4ONDmgLHyEcFiHBblRFXqfNzJAbMrGL6ewRoLS9r/268DaG9
YI4shoUfxcf5/uvylJb4Hvl+5mJfTQeLyljnCLuVxjFrHthYujt3dCT3Fm9WEYd2uOnGvIGDyZTE
R7yb8TQKDZHnsL6kWn8HkAJk+iPauQ6C+GTwtyQdif99KV97YMnocvKmAZDwnOqf1TWhUlBKYgoD
BQTwmy4YT7ANR6pW5lyy9iZxNtENBxKveXCfSMdjG1c5guXz0tGzaxkVLHok0mlNMuXnk/4YoSxH
UPIgcxYXEM8Pkh1sdhQzuZ/ZzscpbI/AQMVStL+funnYiYNrDrNc/jWtzpQot7gz8LLta5aOT8lH
ATJSIN1tGIzQgeylnFwn4K1a3lDNsjpSNTE3UKrptGLkdHoqkvGXgCFoX3u31Vt4ou8+LzAFTZZf
2s5tZFTiHjTaFdWtoM9i/EpoBXUGMGQyLa9JVNQM0spnZqa/Le28OJqkU3GmHCLvR3aBNLHEGSg8
/suzd/MqvsrQM44Cz+6oNWn/TCUeoIWj8rZgaTkWVuEhh1wPrGQs3trZNYGmd7gLEOlFesi6lINy
ASUFajra7fE9ei373iPYQIJ4A/Yqc13VzZGWNcX1lXkQUsgYus65FO2MjjqrBFGyh3qcR1eqUjn6
sHzLKI0PAitN+PiOu9S+F57fiBxu/WOSfONt6gKbkSCeLQ2JDeVwk57QXDwH6Z45T1+yfThfSl+V
apiNCDUBHXg/swRV/6hw1D2Kv6fLvk0ez5Rwg+7rhevbWfR9VxKOfeeYdQDG8L8hbJ63UP/snfy8
xlpC9x6RlbaU6IyU6+FXhDxoZr2onmWsGJD1IvQRu8Ld7gyaqb2flZ7qFA0J6wTcM4eK+oasTo0s
YIC/UwRKUUQ8gFFH4AsMnhpEj+ltmc2t41lx4J0F5S2yYRRybNiL/9kxVg3ChoaCVSdw+xYYWzfL
UKo+3qCQp2tKKb/McUNLBCY64kkwNI/z/6avl3Vo1IhJm1ZsDAoZuBdOJPTRtKyIVfYdgkbZU5xU
6xBLS1Cx0sM14n5L7lxns4ATfWeUrMUmGQP5Rlk2XBmKs66svXxNjP/TNllKHUr7Ya8frSuoFjXH
7UT0ia0erRvR9hb62kMJZBvRyFpVMNGOU4MWPlOwz0Y3KSOSHQhJJMd5NZ/J05xBb8OtjEgfYLgW
E9QfohTZV6UyscJd6AOxdzdSk2kdBRaCsCnD9qyu5HPq4UTmYwngVFIZWSNP6h2kcKh0xYFgMdvf
zinNPup+dCSLKbDTrWf9k+4JafrPYoaiOJuw+QWc2nEmfen/EV836ycjZT4NtgXc3grzCJjibmPD
W2LRNVdPzvGuScpDYuTVsU3uDXhTgOecm9qfOO8YKBIvOfg4cPTQgPHbPR9Y1LGbZ9PskpJQrbh5
QjE99rUvSNinWcRspXNnxB3fHsajlke1jzr/DM/OC5l7ln3qT5IKwOPsSzxVJcR/vVx7rAHayu+o
sfdR/cPTjJJk1j2bs+ocBhG3YyXURGc97lHUcG8Fa1joYkhxVo5peyPLn1VQEnommZcdQWdXVD9t
NQFv4G7ScwqRWXdbZVz+49RbJS1rPGVqsUwpbmTGnZ+KPsuQd4y8MthPfORh68GiY0xgklwaSDyY
HI3OeJuXEFaB2e6dLX1a+XHD6gdxFKJ5U/ls9O2gmDzYomBK32LTk5h+8s2M+wTNhILwrOH1HSFT
wZl3OBQZAiuhAG7DiieuaBuGwfzIYFumYG8oBTGn65fcor7FFP3i5DiZNedMIPcqvzkA2giX6wKB
zLMkZdm3h+ILVIrLTZtTVKAHvkAZDWsvAU7rF8GgJytacpMXvS5bfJMS1VWsdAb4K1w0LTYFejbX
nRHORs0ZhsMfhqFC8ANRq+X3+F4k7C6VN4p4EQ9E6GOqreGUjh/UXPQSss7RxigVJVpvdTbgSnqk
3BwXD2RXUjNQ0jv2DbSIZVaLzP7zmI4VMDyxmTKjhIpsCERknuskxMpnxZUOpdtPnwAYUlu2aA0F
hn59w+OU3BG3LoUrtxLSRIzEkKB2O8K7I8E66+jRUvRTYLAno2m7QdZU0+dN+WVhzggDhs/czMEX
bYG2rQXg7QfCLZd1G3Dd7xBJqLJrNo030490B6xQ/MrDN/mPnSOQVYLLvmQg3P3tI6ZBY6ywlcP9
V/imboAVE6u+ur54ZhQOK9JoWtVLR7sR6i4zye0zYF/AIcRRJvg0O7XxncbJXxEkorX6mZzggeU0
AEzGfd7iqwnkAsz+WsaoBmBg0ZVhAWoK+52xJtEjN0+Sg7ntt4bkpVfCBW5oaz5BmOvd+63toh1S
lpt2STdPq/w6JVW6lwhLeZ84sGwt/GchBTbOhinzh1pch459rC3LFvXYB5XqjXqgb+mBkx6336bm
vmzLbLWJzIx5jNEMQiGJYk+ZvhgIQV5Quc6Gewn39Ytz69LMh1755PHbuvdqcEWgFaR67cG0sE8g
b8tJeJ2EXp73MbSV3JoG+q+88ZMWhqXKCgTKJ0BGHKa69gH+snHQIDylSzL+GNUpAEx7v31fw5ZN
vKTVgNt8mQKIzWNtKdxQ1XGxG2jlS9SOJyoV9fn6hPrACC+czuUnoMADge4v3Bj96eVPUsWI0j96
Wuy5ULJVHm/PZKThi4Gp8yMhUZOaPn1RmWaOicwGDicVSrKA5pMMnnshO+VGHmdgxCuDycm8jbOH
9bqMhUekhSZqhObFAO5x+2MYiKH/XG4sqzgCOMOPOI0XodLsPgVkhkRBdOm2yB63h4DQqYGN0xXL
YbcNO+1EWfaFDhzf1SzVSHHyWspX4BX4dDR7/mXSRBfUl/vglOsLlVKBJqrIYtCLqTjIcnVx05dy
ItRfEJ8X+4Kxa9C/bO2vShQrNaPtCU1qVdBobc11ouNaXjEqpQUhKDQ35qSrUBGSKP5MTZ1ZHjMU
SVMBWH5ZsiuDX7SBNc7qGt5qnRPPM5adPZcsCBZ/iVLJEX0CVbYJlFBjm9hODzNVjKsVqXJr2tKQ
ocwSXYGLy7zVF0XFD8WdBzd3D3gmGbYEUJ4F+UR1x/m1vzGdoMvTdqUVkNtaeWO1hVBaZ9Bc7H3P
vS/ZP9luZP+PRUP6nkCMbTwWvT4Z8w+Ohd0cISiJ3zpydP29kpwyCaae9NZ7aAi9CQLodVVyqKAT
mWbNY1dykTvfaJW38woT8ABGshBLcUZBHLVJ3PAnfd9AgOanH/W73ushxD0ferEUGWsEGApTeJEB
+VnHWTwiCgFG39TFUnRZCTmUWYIqtdNSrCKEM0wFlPArFenFaaV3R17uXU6PH0vx+wcmr5Bv3vum
POrFZ8oLCxfn6LwK/CXRZSSCxrEC3p07GaNsC72w/7xx/i3SEJR5NeBBLDYXSlfJfzMUCAEwtwLK
I1Si4w+z0SsiZjloauyzWrsqVYJp9mtPMBi7OpYUkXgmkH5Cjswu06MDLvCbKdB/0s0Dc3Tv25fx
VzrE6/15INHR9Qbl0CAB1SlfXUZsghJmkTbhchVdZeYL8OsK1KQuKadFKDzEQ2INBob/EMGiqUlS
Cr4KmP3WIur963g0gj1jfrkZGJIiSQlz8wXlf5ysKrmMbyVzPJ0PWqoHR0JIRcJT4kvBS5SOmoSR
KNuPGAD1pnzRCptNUejJyjRbgpkK72ljt5ykx7G5bqdgfURLVkIw4AGIZjFPRITiZqTJ+Txxszl8
PbY9Q1bIXUIuCRGNBV/vo9daPPZo+Q59wqghZcFq51Du384WaNhP8RBTm/quRh+GjzvNjnUfiiwk
98tj6I79oR7gzO62MNoZMrdUrmP4GZZrbG0rMyWHP+eiNmpsORVnx0RAFdjpINMmjvUCHgsaGIyT
x80jwM8ImIIj/pAleBd9w9609tl5GcUiSMcjq9YvYMD8BGxP5MZtEp6rIVgMKuS8wGP/N9NRyNpd
dJHIqp/uK0ru4g45GDZoW9GLb3yEKaA2/Z7ZThvt2rXZhjM66rQfIDwAheVpl8y4iIG1Gyh7CuDH
Uwvn+gVUlUJD9pnSFqTu/cAnzLmsDLZ9cpzj/xVULA4VYRprpWBXqblTCl8MnomH3wOWwWMGv9fc
mZ9n2yzhrfXESvttRaIK/9DRjKR6wRkB+XdhrzeBEqVOuPd9QlJf7dkUrIGIZXIEFQCyOWLfP3rU
8b8mMTKkqcJ5CvtW/IFUFPlJFwEX0xHMbzdgdgcJRa8NyeZDW8bNTTvIL3Fo0kr2VtvlNbox0n61
7OcJZ2S6dBelZnRah5gZLHcDcYFA0Oxf0Bgcl94T8NVSN4wxpINLrGzSXafMzRsh/FCRCOlHk8fS
724GrekBuTa4990CMPcvNK/ZIz/Hxqk/Be7lVEgmmbVriRGa2CCx4YiX18NPjRzBmrlSqEfHLLYD
s9iVlfL8tvVdMbZI9atu6M17m/oEbdavf2joIQSjo3zk3n7wLQFHk2AYG2h0OXVWoxR1DV+7HpuW
5GZdXmMtDTEe5b0L9EHXOvTLVvFis0NsGrlit7vy38MleedE3HamvmCXNTuK1FcXg9J9UyL0/Gqr
i5KkFJdAOv24RgpAIEQMNNh9Ufl/hz5XnFUHagCsDaOqIQy/ngNEQfYbFMOXa9zbV1FJ5LyWnINw
iC6Q2JidGE/q7rl6D6yoQ2+wxmT2o5rJMl2kA99PMFxuY5J8pk1XUHSSlvUaXMIFC+Kjl44LwtA+
jZSnff3xxsNkznLF5O6BogQEmURL7jNyllzxcxGqfZOesGJ7g1ksafYPtCfugZkjmTNSNb0aJm2Q
Z+Bud5r7/16frrXqE4tlGfImNizJkeT3ZpaJOXWuXyHbXGdLSQusr/MHWYWHVyPHV2o4/njmhmya
0kgBpJGae+lSptBEVI92iQpEJt7dq33hfwcCjXFA2lOXgilfQDcc1Zrs49b+7Kzo/zNpMBdXddtP
5yKi93v1jC8S3S2GgBHBnUjuyvp+b1m7o1qpwv6mf20/aGHZ0KTWkY5FZW6325V8FuZG8NkHmgpj
IluruKm+xr21xPkJx1xReHnVdEvsDCxssG4XfiOENlTdUafZTXwxnwNv9FVNm1v1RuxATr8CEOVV
LTOMfSFFrag1/PIjB1YmUxpqLK+1g1RzX0n+nXMKFQytsc+KkLnqp4IKu93/uFvjaGwg1SZEy34S
cwXQL5q/mbiwiUyC5Ubtlo7sN2MngQuZ5kR3crhKowzR3VKfZShNb0XV8WCxeEoOV9lflvDhdxm7
fnT74gwLH75coGYAgKIAbvSq0Vb1x6zvGsHfUZMn1LAJ7tpjGEBTnJzxXIaVA6X19lC5owgg4vKg
/1CVvXsxhKgtvEgcTRAzbdns1d7+rjrJaDBcZynP+WhrBTeIMqDR9Z+HkH+ndq8IN318pG3xzWAp
0RSN5XNHZq2LnVyjs+q6Asq+go/GPRqwEQSGzKTQMrZWceVumykeY55iHahxT0XaiSnuXyaZ/w7Z
Sgdo2IBu3zg63kwj0l5/FcBsfA2HJlU6AuST+JP5O2jRJEDg2r/vKOsBZ9INmWMHnTkfzpqlHaVy
UPnQrNKgGIfZ3NWTh0KDbv1ZvYKDYJ5dcEKgy8j/t7gw1aimTOuopqgp3lg0cxflsqFPz4Kl8Run
nuQ1IRXva8VKRiF+ZOHhyRP2GmCcMjytv+eeZ/4kSLAg6oEJ/SjWIbOjgiGIY9MlWUn0uuFAtlqE
w8WLKH7OtZgU2WAs9JJrc76ob5ec1I6e+XQzfXyAYfVE3EjoZF4krNX4ul7ONh1BxKJjGKELm/Mc
fBQIkZg6aq3zxRDBq8L9BCaz4BJn4BJSSVnjtTadNms7o1nyI74l+cT28vwaimBVBEI1X7UYMLMF
dmNNbw3Ui63XxzncDnrLZ+J88d0Qn0iMIN8sapKMLRtT0l6VRK2mNJbW3viA9FTNpWcXIDbEOfoj
v2+dQjAGTG7ASRrj/SBqBmnZOqBDanJp2AoDecdpywnA8OgfWZOEiv5Eg1IRH5UvdU3kaFAGCOLM
+WurA31J5GGNmehHK2melomlArxVjsaLy1MoZWNYX77bd0MXeanTW8QuvijBNZwSFbfMVY3jgadR
QotqQfTLseInvYI40jeKqJOSDUARC7DUD3sfpozbluknYfPRsYiH56sswXz2IGWubixQJtxRifcq
FrpR5h1D4VjXxpjxRGjwWwpT/eN5oDRK8QpASD66DZ14xbn1kxrtr+lOJXUsxn8F5aA3eN83ZCYb
QVDmD388ftlHfIu4PFL84kMaze2U5CsSjqgI8h4pDLzqWNofHDko2JHBWSRFw7baENuQ6N0/qi0Y
U6gyfAvF0846LQsN7p/uAErh6eOxHuyDEcqqRnvFeO0u4V6lLKOpq7+rNXTYoCd7FAHnHZhvYaD7
jr7LMOlGK3cyUR7gh3LG4Jl8K2tQiwRw8aYtSO1dxPl3LTFn6cqXPEMFSHCAcjnchhUxGTm8rosg
Fuox9xjil6FiTAnhdnAeJQDcyl/E3AB1GvPz3nqm7AWjfvZQn/3SXxXj8MchJcqLDjwIeAzhWSbF
67oegkPZfCFXeUiuRf+d2Y8DPowUxMzvb26YBcPUpBkQOpspLSw4MMGeG22kWrdzx36eLDhasMGM
EDP6eJWq7I/0qAooOJOayMmnaG0CCq4u6boFc3zKVRVOxTwHKhqm4froFoY1ZRdaGFOH03/TNSDk
N6DHKd0ID5NrhfLD7HqLOpzOw+fNxpuSxVA8PMmmRfcwiGaVhVOlJtVfpoNpA5vFcR0JcgUAcuAa
081CjgvYT44H2RhNJzD077S9hxg3BYU60fcUuYEhAuGAfA0VXJUb7MmrGK78FbrFx/m9pKQEK5cq
p2TjGHDvOcUUeLiAIN134bT0A/y5q7HmEjr2cGNmYCbV1wJyauay2sT+OpFALR0iveZJkJDbgkWk
vZjaLImcogwtc4mWRU7EaOG94S2LOE1jpnbyn1kcbRlrjQNf+/sF3KMDJDQfqmHKLj4XNCLHykUN
76E9S26hid5qxRS93KGAxT+f0dN1deoIueWXjv6sEUEH6G9vcw82WJQ4aB94k6SxX/NF4nv6qryA
n0sPbMVNHXsuJ23WIy6tSmCYE/Ypn/Ilr7e7Q8e7mHlrWYJp4ZUuUKpMKMHXabW+dVMceBk0DU2Z
BvZ9J7obVpt7l6Pzw7uzxKNia3RNgtExFbHyjb4IUCBn7FigOjstzbIIUqJep2Q1BfJpSo6x4XCO
bjVHiswL7VHwK9xeH6x8f9Ee6Ftm1flqtJ/LYaGeSr38ENJFeWrUHDo/Jj6ceaGKwbMAqoLWkWvM
EvP+brRCw4pd4D1x0XFC3o5aIDdBloeeeUpgvejw33769GU9O2fF7JNOBJpytA7AeSM6N0l75wZq
VG0j2xp/VcMuE1mziW9+iIPZ9X3BPh+/6F9vpl5vStdZf7mfDcJt8s2Apkth2+mTiTHNPC8gmxgm
lT9kyBXKGuuKcNGzA3oGj2JBsNoiW3UXeOieWA2LREL1siEbdvQKK2j+5ySt0KZdEgsSExB7Rs7l
Wn0ygiBXknVwcu7KUkaRJExbSyQbFEiw9RIuBSJixyMAj9DqHawQvwowI6kGHAWXBRakm6Gw4R6/
ginyPjzmHstNmZODw+CdrJgfhm9CSRugS4jvAmIZ9deHx/WCtQCX9sR1cUFQNoSku8//MBpKBd3/
bpWlmUB3tEQ3xj8wlPcO+tDw9xl8CR62adN5mAFpAvRajuzNfyN81YiECVHIqoC34dGZhTd/tRmn
TJVxbXsiuNhsBd1fnbHkm7bkTlp9xqXexlfuROCi2/db+BETmoHdLkloJhamnXK9sFcK8n+m+xGT
NTi/TdBTjuigfUabuTCjHUO4N5GZSm4SO/WNa40AEtW3sRYxHioJPIfsqRtuLG8WZo7J7BjsefAe
TuLrQFUt8wE0m/sFkqog6blEPc2YAbdaUa4L3eTEGF0HMYcYLCMoA/+uo2KQCZbCChqj8OhTkInA
Nb0qD6DdkxP43pbMiW0iASo0uWOngMeUh3aK3zEEia+UG9Iat/piBlyCBtZgIN/T/oODKM3dngVy
M/XGu3tVPEjW5+lOfiYjRvaXRTZyjsyluxJPabFq/o+sbxquCJKEI0A4UPABQmrZ7AUGeTrLMm9w
ZtKX1rWIfD0f7ulXzQxAx33umnvRfPDxdJVDd0S8ETjn/RDLRuVfxLNiMupT9LHfhc5S9Kq063ea
sQrF3anEwPCWtu2zQq890G707Nhw1iBv29GKVDOKgkbJHyAhGpEYUIywFDjCzK/UjBVWOhq9Xe2a
EIVNI+sYeQUX/6U5SvXBY8Ql7n3tE1Vx9hhkyLOuUCmy0FL3lSynbEkc07j8RcDFU1uhjWWrFRIH
Bhyhp56Ir2cELTddkCRfHYeIp7z+2hNvduWRXnOBT9FL3ZEVzjgD5WsAFJiiSKmOWASgXissmErF
sD+1oxpkTK6fdfyO1++nJ+0tplKsO+FHoFe0U3f2GizffJVs+3wJmrmqwoweMLX8e3S3AUSx2qO7
RlTfZOOoMgPu9xkvNOO8XS2MfM10JwLULtEWtvLqEmNmth4PYuMY5Oai1PAOAEx+XnYVW/x3Q9Iq
TO0fJwx0WFv2guq5xIT29LcziftugE/xRu/Y8jnC9vseVBfklJV3SLA9uGwDl62XQL59QgC3SotK
O8SbNgeZ03fjCR4snfSvlzDOcf/6gr+E9y2/1MW5Adj+BzfsHLC1YuRXA7U+n5oUg2HZKDQcBqMt
TJEF3bC4moXWRrnu7I91srrOITSIxRbxI8LdHJrcStENWAaW20EvekUKVfeg7xyg/lw7FTjsMtGO
GXNmesB8MurCzGVH55FwOsyhdVn6Kukg7vyQNxXtnHx+ePsq+KArp3MxM8kNSArkggUjUpSq/r/8
fa03FTxAtWKMmxnki5gcZUjwHMKb5fsyjZvRFlpA3Ig/fLpeaJgRLxZcb9dtKZ6GJ8Z0aGQsIg+a
+EAD8BLAFwTW0oXzzp7QfmRgTxOAqe81bN5lOzLg83IcBzsDc3RO9QA3S4oCIVVhlgUNggbZs2AX
Bus8w79hOCX2m66DemEB5JuPW81uuFtjc9HHXPoYc04trkJqL+IAHggUTf/DGszerDYQFQmzlr6K
GeToiCLZKQ2rnM5Q4UcT3GRYUw+MwNyXSoDsVbGd+dFhXgPG3b7iHTV/8ixw1ViLsay/3rxAbrwC
i3ffh02YP/nTUAiT1KOqOf9gz1cj1VTffWQJjK2vtmj+O6IKzHdrUbJo3Joxo0IwghICF4IqLjEq
Dyb39tpQp/s8zCHoZqadEYc269Blb/q3SlC/pQBc7zoG7E2//pyKQd8OCFM857lj32kQIg7XA3Dy
dI/mIrhkKMXZNlcrnWFryNDGA/Ux9yclVD4cRG4seAK+wWgr3p5gUxl2cVDvhGZivyR09VDcZagD
5wNpoRz6HOQS7HN0tzebQNutk7/jXciCX1XkgCfJmYY22cWFm/73iBgoCiHW7h97MIqGjt5dEaOw
SY2DkKx3TdhzTDgccjxtToWtd9lwZwyLXnC+6lB1lCD3dR270UK1kPeG6D4sEuakQ6R8FLVnHFd0
S4JV4TUCRRrf2v55MN8UszsqF1KmQ06FnjBu4ZHGtyBLslmmWpPwxadN1pR4yRwqWbP+CSK8KDVs
TMb8C8a1rJXSqLJ8dISOKy6v0O0Oq5Zvrc0ubEyjytcOcfXEp/7o406nFlrovEYAzmVyl+Oh21IZ
C3ysKP67nPoQL9tIuUbyPXOw2Ww7bafvjv/BjW/a9TT1tkLA/IEFlY+fBCpxF8KyOe1lJb47qmcF
XWg60RrXAs+SyfBF6TcT0EzgJ8+cOkT/Hkbh88zEPKo5+eQEojfBem8L0h6aPH02C9f5QMQLMZe5
Tzm2ZHHxmM0DsgZDXtYKSDFxZ4Y04RW0Tu5l+eHxkpCRmZzDvggBAPGydKcJyoxPtZJz5Vg+dl3V
3SyuaPwoKdJES2e5LW2SAwUHo2wHDI9PiQWMpbmBeyGZfSGVptKzJ8WKN/OKSXEkkexjYJ3fsGz5
E23k/yV2O6PDcCfa9iPQw3skfg/ICnFoujZ+VusLhB9lW9/XqmP5KbYfQlu3SzX5rtD05Z9296+O
7LwqEtcmoQhEcjjZmm2KlKymROtoqYBq8+RynLrBD29S3bWCP90VGWhp3MT6Naj5tgdV2BLsNIYZ
dpq9k6/VsTPpkfVi5zP3DRPv0hyIdDUGmNhShO+p5QJ/hqsUpP/y4cRbjQBlbSgoGLWN1hLLcOjW
fytAQ4cvcPiJVSKDgg5KYXABtGuYapZS2IdN7Je9UcNaF/4GlEFkP8oIZ7/YtqApgdVmsVITaPR0
jgY3WTStSK1s+BgU3I2GDjM3sah5xywcItSctsoGsOn9Uo5F193XWWp/xZZdnyREoNsMuwAjHl0+
9aFQshgFiBTwWdM0PfmcXpjjVnw4R27U60owOHSrKI39Pwz+Mx1I2zqFMNiANo9HDN/J9p+3R/Iu
k/Q+7x19r3mqX8I8U7k2fBrf2wRkVlw6zqypKKinJkXrJgdrt55qZzbqrgj9igsZpUHz7+At2417
6dJsl4n9W5Pqh9wZMtuM/2/biMJHjBw0Y7UM3ZGIY4Dw1Cp9ID+40mOALmYhX6YdTgvTKXvJoapk
CgUdad1bGzqe79ORlGXFDjs36guhVItuXxwrGSISAB+wFNX3Q2qF9fZTGmEZTC0qKqNOnyWGJ0ik
xKwd42L3XeCk3rVb/8xRkBafqX4tjuv7CdsVC7+3RCd/dXrzrzRDE+iMhzkxJw5HHRVzXIMf2UBU
+MH86tdfjZHFcUu0VLutAOzt51WILD7TguGsYuGokTNi/pqtfy2/vnaipx2gGzSzlKFWcoshoL5e
Cw6XBddTxLenCJdNys5qNGCxqobJUF13Ji/hi1/KgiGfzG4gu+DCRTAdtFo+n09vAo/XgCSwQ2Is
OA95fD/cOh53xJOnqpJiPqxBMC1ps8v4qHK1LvVxvTu64c9j9puXHuLIaNXct6i/GfDstHl/2zbX
OQIKyRrz2k8DN8WIS9xZyKwPth/lt1kibj17F8/Mq/4w4RqB2LnFFUQQZp2qJeJhW71Ga7wMqH7G
0g27by+++bMut/ORvctspbLuyUAbQbXVc7ek5vY9CgyWWYtdYaPd7ytESsmIpxdKbwUAB9mII0o8
nAE1ci1HlYqfvOGnxZig6E7jje1rsG0Nq57yOK9Y8tMgkUzUWJK4pWZe2fXf2FPXrnRL28tBQ9kz
7wPNASkSCvldaB7jaEJF68yVBW1fJF87MeJRsPmOuLu238wIVDs9Cl+d9gGpDUM5/SmE6kmvQTVg
DUzis5WEw4S4K1521A1TCbZiUnNO9E6hqKegq84rlJ8tqN8E+R1nVsLsKCDkrPIah+DMdgPv1nGC
a5DO8r+WxkYwQsBb8ajHe/eLiT3NB8pHEbcie81sqpYtv/ljcbNnWxWaft1pWlLrDdrj8tmvYTDP
HpSit8Ix76//z4HNJROnZyvwIo56EOSOCECuYlcI4nggz/lm9xzw09n57pXTb+K3IekWy9a9v5h9
3CJkl2wLJUJxkQeCvstvlpC4n3KlxLpjVIHZ8O2Wgzf+H7Cx/x4Gfwd546ADBqaEXKlgDeF7jv0A
GmefAoOP2HcL/ISC4gOO473QxSXS2rNwdUEqAArw8zOY570N0GvVI2eugYqK0QRpu9BnXIAFES3R
3JdbJwz55bAe1A76LMuAeIPeKJCrvwDeXtXuxfOB4RECx7SLkEJPSfRVaXs6nPB1cOTnJ+jy0TwH
kOlLohidFJVDTRVDaLywd+CvgOdQtxTeXM3RCbxk7/perGq4onlvr0VtRywI7tW71NjSsrswjkld
d2YLLZ3gydFgUHA/ChleGD4vQy/boWUHJzguUGpm6Sy/5J4WNtXa5lCL5qYKso0qAa8+KEpVR+vK
5+7wO5PKWRpdXILrDNFD2zIyhBdfXqRdUFjYhgCQd4IL3xLdxX1njK19JziolPhr279KBnixROOE
lxb5qwJr11XdPA7qcEcO6G7KY3mhsa5a4/BjgiZY2ZgV7L+Gh5NCNeU+q1xKB2wQR2HBl14J8sAy
8T74vstBjpVdocsJATlsCAX1O/JV/V+SNn2HFRCSp4mS+MNiWpi9/xl3tXQpW8v2bBNR74HTmKCC
RMw+AZ3QRHeIqFIcoCaP83SbiIRYwnp3Y9KOZrMrFnD6Tu2zqzrBhwWLh2FyaieCgCqaGw6kO3FR
MDx+y4NA80gs47D1jUxbOd3gcqcipYQT/mg5WLKFD7OvDJXx8UEfnFZFBDVVX0MvUh9D8cMELnhM
zhHmJHNo00hXLVQqIKzs49/3HekO0u9+ui2laEWbT6ZK6I9XlNPSHpgESDSpbw+fDA+Qse1XKHIh
DhHLmLn2cAf+yVMLgKtvvFQqKZ7P7/gzSG7IMkbryn5VZnY46Xt+1Ssn3uhdEMlRyidntsY1x3R/
mxmWNDcIJ0H/sawHPS0uuU3+mZ1wgX8S8zS8RFn7TtuCZDh5kr2ICSOgYSj72TLyZFK1ly2/Tn2p
fXU00BdvikSb4gABprHy8dA/DO7F8Lqd73WxgdHb3mcwhaga676GBGIJp22tyhQ9EnUCW8fr/JR9
eVTh3f73dD2+bt+3VEH/7pODSooBIMWaRjQzbx9DUhm1zBpIU8K/7Trs4tM9d6OMZBNPisOTrhY/
+aYf3cz6lW5GVhZSQ+XzOnrdR+MTaCEQD49xhj+LF2qQ5ykEQtYuo0RWmdvjFjRGqyhAF7SwOYck
DnaBMLLTqdsR29JruE6Daw/r7sXFz7ShK9qg0CI5nzEK53j2W0Lws1zklunO5RJFHvF6OMjmNu99
SJC7bcsoxQsHprKoI7nSPgidi/7569gObyefDrQpMi137kz4CcbIPdIYYqbfqul8CjOars2KlUJr
jwCL2t4zEK3vpQp2qSjyBKUqa802+ahn5dt7h/u19ryPTDaSGllfnpWBYSqH0ZkfQrgJDp5Gg+t+
FEecbj04qmbVsAseiAdWKUaAPyMN9f9au5xf5FcYI7E9lL+S+Ysts39FW/b7bls9n2QeyensyXAH
TE2TvrIb4MxOFpQ4spouHxJh0BtS+uSxyehBLvKmU0WJBz7oboRo6BO0QAhwb9aZMXD3tWaHZPv3
rhTTAtOGHJWXVN1xipJTGykh1wEaru/SWe0mh8swb9VODqaUql2nBWRhp/x2mqNjYhDXHiLazZvt
f4fLbtZqngF8GaKwI8n30LVKpYMI0NHfLcLKfghDvr6d2AKdl9A0jck3HjiTmXEZSUct7URwejNe
web29EQrjCWcblJopEDcqt/ExegeyRL5jNNPojRc9sTFqUcl17EL5PU6l3R5q6HhXz8pOHnZrKEO
aicWomz4PWVKWlmlWe3LHn7t2LuCtflx6G/roh8t728Rdy7Dkw10Z2vKq0Wd3MvaSWefddD0IQ2M
DqdbC58CO/38vBbt7BPj0Dg41jAj1S3LWlGA6rPqO2yp6tMY5+W5ztGpyUG4OhuYAfRCyERFYawk
sDnyKa9e8EbPS9ZFujT82hQON6ymBd11hcAGX+8xhXzWvidTkv+dt0DYygeuPF8uO0FSrMeQ6O6M
K1HnzSMdq/GY+mQPi6QTb90jJEPYzeaB058i2+crt0RG4JhkHLsB2IIKrcV2E0MR3X6YNBdtg4W3
r7CO4MsOoTpdyAvmpmiSs8EPY0ZvAmcDWl+eXExZUwzNhr9FDJyaW4NmYcgcky5boQI9nIz1ikpo
MzBCskQUYkRjIddvPk8MpKVJ1T9FMAhUOg/tnVsu6qzm3ffS2sa9B3ghcZvcGsSTpvqUVAPK34F8
IwjuV2jDoMQQJfPONacJXpL/lwlIhMyUfC5dVK2wPlG2Z9uJxgx613+RORsFT6TUyvhL5gyO5lYT
e+9xppeS/YVc9tpR7TYQOy9v6bt1ynLWEms4tTUnbcNOL7trdsJv43nf6ZF8KFwOtluC1feTS1M4
R8JG9BpCPQLcusYyUxR0ocrD2oNzb76YDYruh66GzfuS9E+elnU9LkRzql1S+bkLRDaQNNewfKt8
c2MDWQv2rSgy+bAk7NW3Zlnz8WigA1Hnhb0db9P/8KjUPcLljZfmXeVC0a1BGF56lm41kGOtEGsW
sLzJwioLYo7f8GFZzqP4UkCeMdQ+jl4sEHTSmOHsq0LVqf8uXWFLXNe7ggFdrhr2nF/P7HI3M1LL
B76rScK26jsIdfmpdIy74CyWGMtKMNoI1JMwnIvScQBKOj+fLgU4cgf6pv/CEFEosMUQuDM818Yj
N+11eezcW5xImeWmDyZBFjDaG/pU5sP31PQQXi5AqHq+qC3bq2qXqCOIj/xuIHLKNucDuAz/KJ25
hG6uRzLgT5+y5vyN1YfA1J06rFNBqMUGZAK4mBC+CxfekHBkUwgRXBZjZTf5DAA8wPpPNriy70a3
pFLn7ivinchaPat1uCkKkDm7Gw93RY2Y79QDibrszX4TXecvgcYf7WlCO9FkQy4UGRxFXbrE/RwO
MPAXM3n64GiISa+pvDPzC/v+DMgBojXlYpE1p3xDPliGGpwMKfqLSb35IBZ6WalHrtBE9IUqInJI
k7nnLHWUVwxN6LQe+F7ThfnHXwIfTDPzMz4tXygddOaRxkJtQhmKAlpo6GBPJeMd+vxNiiwlTsdJ
iRqsQwAPX/qvGZK2tDI/a2PONAImd/RQkbj5nafgsY+ikoISP/1rFYX3qQ32dL2k1JsWleZW0YVN
RVhAdDYv9BU7+zuh95kALtIlZSRn5kLNxle+pqmijf+0u7JnRbW/zbQV/K98T0vvYGmz2ttuIeAT
kuRCp/sfLQJw2f28NgabTaNAXmRKOX5Lu33lG38Vczi8911OuHIePq6dsAgtDBFWrvIiVNWKzSaw
ThRBikFF6g1yJDp1i0XGIHzPDvj9uiIxNoyES57AdUQgu1Quzoqmc0w4cudp42WBQORKnedv+HlC
Qb76xmb2Oqdz6rR+BY6WvPpzdPDdZyDDbfSH95rWauuXMFid3Col5fmBuehydJfsKfv4zX6F4Ysr
PgHNObhq8X6Ngqi4VyfnJ9wa1B4n3ooN/49+cA8Y0UZOZEUBa81LMyOlIjSTGctMOaLp36wtgHXR
zb/TtIqrtXLI+W8Za+gpQe2EBd7xitAXAQHEnqE6qqUlO56nMDMkLNrW+ipcyiuXV5oXygmrO7EE
AICkQYILNO9hVC6yaqmnqrqGnq1xtg7UCKIlRcXRodlYOVnzaRULqN7SCil/tuWmAoCsQgQbLc7F
HVS7rv0kedCOAkrY9iwmmBi/A93nCJnKs/PiAJhueb3Kz56TqHADEpE2DV+nq9eejLvTwB+/HFwW
NQbpO8225+AM1zHmgmpRzBESkK7y7ncoU5KH/Sp9ldqYnlLWPnNvsaTkuhAAbhGc+W/x5Fsxstri
gcdr8JN7MlDUhOCvGi2jl6hGoZ4e7x/aP379uzHCUf4O073HTIs9P9W75yizybUy2d6IcHA4luCn
12lcB7bi4AjNsWdChb2srZ5KX7OOEVXezz+zO3Rh6aSmD4QU33pgkuv3nW+TGeP3A0E1sZMAbbAw
BAJb/Hw8Zp2ayzjI4VXO3kQKZ0jLHkVFNgosqgfWyaQ1fs9JQKLZFojuKgNCStroaCIEpZyNjAQh
hyvFvrpkZEkezKjU3si/cXFSwFrgdqa365CHDXOtNzQY5GKfPYD3VKZdGBPNZAN4MThiOLTg5npz
t6llMHbTGoHbS3O493WP+Vf56DrohG0213CLIjA3lKJpy8X8qT+/mG+2R/HSYiHR8EwhaEcyCRSN
nI8814vj6/leTgVGTpHl58/N8vsMr+yDgWVMnGYgNrELEnRSPBOKFhOvyMeVhFdz2MtNT1O6M2Sx
h7+FeYpNJNFA8/xUCAfPCJcoS2h9QHS7PX1UrQKlhZOlyx5a2bn9uqvKrel2NoNa9sb/01o3Q8Ss
HFVrOtO5XhrmZgTQV/d9Uk3o5nKixopMordJjwUPXKRwimL6Us5Kz5EymWXm8lMGFm1912Xnuc8V
1chYB0+xaH6xNLvTH1xRrvszCvDynTtsvrP7+9cV0FLOy6O0jv/2XodBE/CWwvhQPW5laYQmY+8s
u0gcBxeWaQ0RABeicgtZEPNsEE1i1vnQV1bRLXaLHu/V7klnw6RXVDWjGZEFf4EbpjEiyJEepQd4
HcpM2vPDkaV3SnP3hlbyA+nWJfQbXKiI+3p+mPlU/n9gu/GFjgyps3vtxjjwGMZgMMm5YbwN3FFb
J0qtETbuH2OyUHZCgxZzQ7a9of7OttIUaeqSSe1trvUa6OSQdGkvxy3XsED/hpoHCUG9/zW2+faW
e+qo6bsN5Uv0x/kqNcZL3H+jcB0LyDiEZVWvgE4K2Z8uGjJ/jphcnguVDXPrdZBIowTk10Oivhqk
rYMLcx0vBGQFlGWEJKmImpXg6r7eSrp9daXVgScLy/GV4IUCfiZuzplvyUJmDV90Jnbkuk2/Qx4m
nDc0PVNqJKhph6WzlXAea1HjSzDg0JmYEkGOLXwIkGFcnn9jA+9SxW85+hnZGwRpu3sVC2qtpF+/
YT9o7OHdYxMx8FPMNAdnd0MYKr1f/22obdYcDSF9hvEysJjGibabBJl9VYVjAtvSmOiWIZma91o7
k0g+UAtKbcxjxzxk2QcruPwLxj0J3ZBM57A8aPaCGW0c8J7PVF7PRGSwbTiK0U59BxXKtqr5s16G
EQ3GXyGS+nuABdIjZrcwwL2XmpGeCxESL+hwplFCYMARj6K4ZEcURf8tZ8oUK9wt3kgbjarchJUm
7GL2ZiNu0sGTXsYFE8Fi/56g+k9F0FrmQ+lILa8fHNVi4Jk6yOGxnRFrVGUsn2RQLOOzlPEIHLJG
dwGOCeOhdJlmn2UsBJI1SHgc4V+xmVJcWS6UVxeYDHhqdmTgWJYPgtJnR9gPpsIra05ZzJAf6N5m
lTllE6aUZxDbmBQ1AaLVnz4CwlJnMJtIp0AAZiXy9yrBVdqzRkRW8GIV8feAWzIhBqNfGcqFGq27
VrolECOPCjBX0iH721Jmo0Bjg7wssHrv97m8NmaCdJq2x9dnQw6P2KeHdpsALM5YMlkezzPyFPNj
VHaiMI9J/C1wnFOgwLfm0aGZs/STIEoTMfQObhBJdXwXgHET3W954e24BnfV5Rx5BdCOyvaHwbIb
Mj0r2h0UEGBJtikzJ28/KNZ+zrwnbX80vhU8nILTNHvWz1ZRCctCUqBZg1qwNpIM4Mr/X1ecfl0d
VcM+vBhAf+sLTGrrezYFtwBaSTA70liurH2mx7yMir3m5XjstyKGpCHfidbqF9BY+mg1vK/yoVdW
r5qp69RQF4zjddsLPU1ydyC9fN+PNF+5yorCe3V4YRk3uG2p2l4ciBEampMb/5LIP8zeQm2LXjve
Cxjd0k3YOifT2zy8jTx77dssNrWIdC4zLygL/PHW8s4oBuSCphtEJQuTZNmjJ+JVIJvytLKx4wXL
nt63okVfdgdHf7yZCiMbBlpH2OdiU+GNeO+tUVZsVZLmnCZf8jd0RwH8V6vgbn7sxoMphjCf8pF2
mo48yt90vZvuSXYwua7TC6KFJPvNY5SsIeElbPMU00uFDNurgHbvYefw9d55fNAL9NtaDxzRbKyK
DhtPmddbX8AN93Tsg6I4cwXEvhuTHhYuCe1SNqAIeRnpEK6dESwM76btff7zMTgql8/07JKW+FgH
ZnFAMYPzPMCBKLvXIqZ2rlyTjNoKYEs6iORO4V3ICDAfI02PxDIf2w0iRDm2fZvbLHuVCs850Nma
0rceWg+ZyYi0NQ1SJD3+blNsAh/TTjw9JxQ6MkJTKLmu1AbdjgJOFQRzxJi3/dWCRBCNncbEg256
fmm1l+wCGSVmbu6HZtzmAss44jQC2rsQH1hYh5UQtL0Ga3xwbZD5JjXgOshG6kNMy9iAD0//izQX
EJ8ydjBBwJkejKqe61AidjqvxGlcXxQvby5y06zCmX2pv/3USnOHxMDUT0LLwxSgbbChfvg9i6Ne
ieUD7VBXjmbENFXlPtQUT4GwjTugGb8kXn+Wjroq/ucLflqzofjiwYZDurmG2oM0DlfoghsfJBD6
G/VMc6xGnFWR1ZZJQ4YUdfWWTMxRLA0bTlmZOihwfAIyiSOPJmAEPRryBBj1414xxH9OEYf+QcT4
cHctxXICdbMaSKEHHBDW5mEfkcLarFPjEPjEfhn48aNlPfpqNWQKe4uzpJ1YLbszM3Gvg5/pdf1M
9CnyaXcgoyyOK21EcwXSC38pwtATFErt/TFhrhpEr2KWBAMudVcU3Dv5TW3QW/M/omHaahyi3wGy
ZoJOsstD89XCeNKuQJHzfXOtJyWSZfG6oj6ldZ8Z33Lg73zhBdHdWLaBdStn6XX8kRDf4KyFLyqv
EuUthXGwZUqFCnabOm7wQBPyIWbiStsQ9L9tZJZrBT+d6S7UuVl8FDJ+W9pfWhfLM3Lxwv8GiPi/
7cnb86O481o3Aegb0ZfSslnnImlroRFerIhamqlL+otGf/8yM63/decrHfZLSA8L11EZWyXio/ID
n2sYZ2BSdtMJJKCe3viRx+qJlPHvZ3kkPJct1k5StFow9k22cOCiyUm7s/x73RZuvWYU0X/HjdJq
/j9nybVceoRVzNQ5W4LbN5TbsarChRlP7HlLWd6cgA4Nag0BchhGc/JdBk+NOY5QU8F4VvWrds75
L7eAYTaGFFIH8ln0NBzTdoK9DdwYxH28K4Vv+3ed2RceLNJJVIyixggpHBlfXQpgWe+gG65wN5IE
4PZldQEpn7UCbM6Zht9DPM1i7ZU9bdRWgk/rIL9qGFpmZRe7QG5EPCZjCFdIXcAYOq8OX66dcGwi
TW36FHDFiPsItPCkEbrqQH9rLlZ916kto1im0JuKdNr6M34VKqMaBfudNoWR4Ejyek+JxTqNDg4P
nz9X73fRWQw6z8Qa/flDxo2Gj7UUkYu7iEBWWsZZrRqVDjOJ02ktkwupPcHocHa2T2+OU7p1m5Om
kPpAOeRGmcrvoKd+6lEFaEFOV59L+M6Wu8wdfOH8Ma1oKcsBiZv+Js6YquDChqxHB7X9seGUJ4bd
EsmPvdYQpJAFtHVmsAYegT1/P7PzEmXdfwJzpT11woel2Oaqgr+VbHMcXOxTOfote+a2dAHeh3SX
NKZy0YlE1b9ikjAK8hrbHsZr+koCtTAfKIIfoAfi4v3NXSj8Oaxh237aSrb9GddS05fMMozUfjNR
IovuwVCA40gP9oYECIj0OfcfEQwjlb1+4tqk1H3+jemDv6qUvbHPLrwY0fvlJV+6jK39sBj+wwTt
BbOAa2sfBXmz8Yiib8jH8N0DUzN5U3/iMTjwSkvVm2VRBHiFgKbvVRD3KlrtXH/xq/n3gBwc4QVr
C3S3g63Kgum+5/+oKIcbRp1LaQRm1D4OZO+U8u1lNctOqqCcEo9/CmXeFgYP1e5U1lHWZ7hPi0tf
YDBfFqWzilR04xFPwr9igCWODvPlVhsXvgQ/NhigWisTbQrsYHrCFf+MA0EgKg1CPreoU9Lx1DjQ
BF8edB0PMjSuQAc3lF8XMUM/Epxfq6oqS4+UukKMRw+srNscfTMRarypasg/xEJW6gyR5RjTmSzE
cXjDuqn1k3Hj7BeHVcc9aIB0aWP819jXDx97FmeXkXnIl7zN8LX9asDbhV5scb5KGRGnnrR9OiTr
5IHmzf4mlRWEORSrG1h6SHVigv/EtQXMgcss0AKE6YaeW1LRBdeQWHexAfi0GKNpkv28sCYUAOPZ
zOWtYHfzVYp2/Q1KQdfKzRqagJHrqxTkJnVXdU/ogchf1UZj1WzSTlceOlXQfqOZ3YuQv6jhP7F/
uzQnS7EcEqts6k+h+lwH2I8hYzG6hrJHK5Kr5yYC/FuOzLUKwKnI0o0j3V5rlkexDoNQC8OOixCP
96kuUKeQA0wtIJvQzqj+4sFdnIrtGbpRd+0lV0Rk3u7m//S+y+bhVk4UK7yv0SLd8hi/n8TCt7X+
ZlJXRwkcjeBkKk5SfD394kJZwV9EBCF3AY676Yf0q/vtKPVjXNvN8L9QRoTDExmmEtN52HkV4CXS
Ckt3r2u02o4gS9mILm9+aozQuvEbU2uGNHJOmQldN0V5sCpXcHcWAu87A+loZY9UoF/DQ/Yt1dHK
YCRtylNIxAfiOl9uVkz7XMzlROdbQzYLVFwZXxpcxxs1b7E3T3Ql2xIKFQ3tD/fMZFmA0gXoCbE8
2ebFj28Q1dYE8Ka+b6Yly6q1J4TbGIU8Pn7hpy0MBnVIdJBIsU3+TDJtuMFd52ISNMpSkVAap6E9
0YzHNKpoZxXPX7W1sFQmEEVgeXyXWQUF63CqiTWkCRMmEPJ3jWF6QTP+v9twrtZe+1gIg5rFMKvR
oKdpMGf0fEPsptL/MzI0WfyM/fmcnvYzfv6+kGOo34/73nZBK3CLrr6tSEYNlUuY2JZw2dFrjbEe
+aUCUOGffB2Zev8KcCkqXdDo6YX7d5mn90aOiECf0bxfhTOZq46isV2j2nzAF/+5VAHpdgXqqfRJ
gP8rdVuw3ejaUNGjH5zInYtfD/udDab9mY7r1qhLwT5W/Ko84vbrukSkUBW/GIUclOz9YtBBq+U7
9ptW2iQHL1v/W+ODT312EIWLA+vmF6lQqzueUk8IT7O2NE3C2reiqvD8GLQ6CaAfspiD6RMiAz8N
P7XfKFar034dLcr4srMNoazc1CfVGouGdyvBzrCKzMO1PCaIUE5uQXjFWlkV14ASgSm9hxxT8PVH
v3Ek4uSFTpJEvr5AgC0NFZFGIFH3YeZRCkPZviIGlitHQNMKTlkI5IueSVu/LfiB21rz+OtIyE+w
e/Eb1rHUi1RVrh5eAzy17lKwMXj3fn0lWZKPkUWU0HgC47lL4h+8lLgNFjUVG8hwlkIHMoF1iDHu
s6y8gzehuEI+rPrYdw7TMIfidxRD/LZKndgvxGAgcsosxPzExsyA9QtSmtLgZSuhbquI0BBlnkmS
IPaGaGQH2aB9MY4dQ7aRWI3oOmLArxEAynLU+cgtTlqOp3lHl94j2mli+u7uNnknQ82lt4hMxGAC
YpTXfZb6n1iWPTFPZkkv9QJ9WFNaPVBMURECkDYuAD0yBI9pvPip31Cc+oh7UrKJfpLVIRO5TGJw
B23u+NX/KM+xB+76LyOPRxY7c+stX63HleXxDwnUiA51A5joZG5wAdpiiCc49O9eB4704rFC8suX
0VdEDQhfDU7mtEflNcBW7ptD9jzWOTPtn9wRLv3kTfJjEjmq7LTRr5ulFBAJkJhV32elhuNoRIzV
PhgapWp+WApFDqmD3FVGo+T0Gqn+uzbPlQcvas5touY5s3Y++HWTurGf8WNDrVMl+YaX3mHoX4nT
dcY/fBcCXWtoBKZU9P2WpTm2uqHOQhm+2cMIle99wPnIYoRmsRixfi/riCVfqwB9l2pOOeTPfS6b
hxwWeFn46rXA8wl9gGhQtBIAcVVvK/tPC+PWuoNLo3vku3/pai25khKDUcmQ6RepEb5Tu9WEv1P5
jaDgd3P7HL6O0wfekASmwXzQPA/0xXSGKnyIb1/UHs5A9TRibd0qyqgRTCTfKeDGdw4uZCa7xRJg
AgxBVSSYaV6ObEDtLVS9ePbNRYeq2eUqObqt1Y3ogSyj8PcPaDUK9y48EzTU2LEagI4NjIYWmc/K
2ozPNZOsxlmc/HQKGEfFZ9qL0bO8A8RZyAJj6t3hSUNl7v/JWRjl2WbFgysuDhjJZEf4VVzYwEZj
2Sby2OtAcFxJ2wKC/pOVqbXLi2Vs7eDceBziI1XFrjkhBNXd6DQUAvZC+BbbdWADZYL6H/g31VDw
UqYM3nMmPMTviNgk5H+36uYu8R4c08qkP+VMlh/GtUhx0dTGSQ9TbuYu4QB7DFWQTW5WXqIIvFty
D1O84hVksOaCja0jR9lZPTC1btkgmOz/NAShJBt2MaWsuhJ8yIQOJrcvwmHEETAJLSOlD00eqejj
s/pTuqnVBf2CTxBPJc2vb6vhe3JXoect3QSNIoP2pNMyw/ZGYmQkRWYEzsrFeX28cr0nNtwyEgL4
ReoLlJYMj1G4qONV4YPhsF1IBOf/wSDkKL2Ao0BHgxvj4lLhee+Ik4ALMCwtt0fEfkVkWQG4Pfgk
3d9jOsFFgAOFOSIUv4ZmYCVZW0KqPFBAPKHfpoU3jaO7jH/v/YKKANxBzUHMeGD3bgOgj/NrLrYm
iY8PCoSU78WFmPRWACG+veM9kmClA609MTZ6HSVaM+TKrJeJhoOQqt3Rk7kl4Jahf/zPUbwIKVxX
aZ8/hC9n9T6NwH+7FsUVSjpK8REHRmt74NEQ3ZgezT6gaNiiojQovGdQy+ILbu0WgW+wDCWFkGOk
EVjG5/0AlBjQ8s0p4fACZ1X7i8+MmEx/dlHY+NxPCte4aGnFd9wC3fXVQgQ/GdSF8k7FOadDtFjb
nDNJAXaiouyABjIuWS45bHIlRbVMck+wIrLQDxhA2GFc3gXFpD//QyTa5IcMVk+V+GPxwOhC3hTK
z8vcrBeXUWl5DNvTFsc23VQS0rXpKflCUQc5rzIqTAm6E5Jeo8VKf2CfyAioLXnSU088e6WNvSKl
QTSbugmkMCVs5n5v3z8x3sA76B0FgbjtR4S+JWKHPTlc50rGZTSesFsRwlbftNxNtPD1Mgtiil7b
CGHtfxJ/0LbCnGL59iHhQ2Jl3P42lyNAvluY3wKxRNgq15/VrAwu093nbl6JKrc5mFg515yk7HeI
Hlsj1ejhBscYosTDGsF8CL/2kGqnkv1hzFX12zfzXhmuHpEY8GbUqrdzi0mXh9P46Bxd92495KFP
WDHhT9rlJD23i0PLNH03MugLrP0lmYzgSALjfdCMWqo+Rz7L7dXjYWlniq5nsbRKMnFhWycdhsDH
MyllyI+taKRMP0W3fqPR5KundTlOR7VTR5uZI+q/TnjsR1/LTJ1AiSkEd8fpOsjWVRVjS+LGk4IE
lla+nGSReDVmPPBGPxugvLP6nmBQ4UGPIurD324x5+n4beBOSYUQhHEg2aHKdXEgrOJ9j7EOI76Q
ezSoBwzSdIXEo0JR4EpHqtgbjpe0WDqcsU1RJ2UzJLzEiIRcdSyGblqcXdYLPC0ktiXiucGniyGB
yoD+5eOicJWrFgDosR5IPpVdfeCeKoyODBYDl3Yc2QK6f1oma8H2KBdQ/yr3xuGd6irvhn7vNfOE
6bFOvCqjZVkpwGXAx3G0KmmzJID76ZkypOU89LPfLZ+DKPvZUE+Mc0QS0R4n3NH9BuUnu88S5wcg
3zeiHLC+1EOfIxtxVj1e9mUwYXPzNny6Q57mjXsphhVB4rpGR+ew8EFFen4Um6HC6RIYuD2r1tv6
mjjzh8ZLXT5RBbXu9T7l9pLnpGezDVpdsAeYku3VlXGtLLlE6NS9ApU57nOVqY/mJHnxN2vZ4ZS+
8rCJz1MeHLkS97SuELU9lPcteaaIJqlPxb1tOSq8Mpuxx0KRRxBcOjD95LHgmguDqakEP+m7KhpG
Z2p0BKbS4w9YCgvmWGPem0bMdZ2PhWE8I9qDTJsKoJfMeWJIyc6jUIPX6/eD6zbno6sRuaxCXv8B
l8tnchSc/z5J0y5O1GHlg+o+BOq/zg3Jk1ccdwOn76ZjPr5vi8tWW8HnnRhFOSvKqDKmldTiaiaV
0bdZ5wHhvbZtmrDyq+cVGHPC2uqjfKBMZxMfMS7ZFE8Jn41HIjtNsAXWE4b5emRfr8Q6wcdy12CE
1VUJTh1jquvn9fAiuHPSYgkiMFS+xC6wJZL7GWA7W6u/O5LTb0q8v5dU+i584AtHkBjxcZ/zfKdp
uU4D6NzNuExaw+D9alw4l4zWV3V4kZiL+j7NeR8ZClbkDmod/1G6mTyskKDa8s1cPWJyB8cbThHj
rY2ttsFNLtP7rpIFocX1mDax5EhfBcXwkzH2zYQoCAKcdCrVI/XyHvSTTXbdG45Q9unZ44zRW3Dp
/LKYwX1u4FP6YmfY2/yTlKqppgVoW713wMB3t0snTCvIS6RkgYIjlPdEuCJagQxbrYcfB33P3izn
JTUWga34WRxtVm+6eDm5lDdR4RgNHCjOH4brdF2kyWlihg50TXRIvmFA93uGSj+FtqO7dKw9R0Ag
rRlpvpuxVko0O9+NdhuPR4UDTwzlSXrsTlwUMMfKy0furiwDIVz0M+L449L7iZRDsHnRpjAs4Hzp
Jp9f1yGV3tXUX/dEUArCPIVd8+YsxS7mk2aNFnv/NvX9sMJmnJY7/NjveZjBmKPUBhKgUYJLTth+
V3UFJcezTTiXN3HNaS2FibnY6eOTNLhghveYqKJitxjIpLPG5XRBH/Mcl4bxA7/q3nMDyUaumbRj
buSbdPMeMnM6orxy5/oYod/G2WbOrVOqXPigEO6iCPoSADFb5VgmwisAOM2p6nAs5pwe4S3BjDpn
JE7aShSE22PPoU0qTIZyEYdcQ4CTA+fGCYUlwyTg/jdZv8eBCQpeV5pekKuIoySsGwCrstWt6pDY
XxOlAQLKZZxYBU7UHjh3HBJPsIoLqDOp6UCblbdpVp9sBe7bNdtDgiAlZonpLIlCKqLyk7CYb6LR
e75/gVFygYJ9FN6WlUULZNlWqb7Y2X361sW6UWeWcuvhc9+AN0xqx0Ff8WS5gXgN8COsOPbE1itq
GBaC6I+HMur4RMt21uzM0pf+Z+7smkkWIasK9H+Ej06ZpKth7MIHTdmAevNYpmSl51H6Eq0IPGC9
sdf14e0CjSnuS8mEyj61kDBvLnbesdLDcMRMA/tFWnGIsVyVaUqbnCxzCc9F7YnuZWu2FdyAemiR
FnvK7iaOwEFTVH75O0VWBdmF+yNFA6v095xN9/BRF5hQuCaPMbPaj4efI12Q0B8ZJBh1JE3EonF5
O8hDmkVqIDfs1C3hGxOSFFmBBLpOJCRikGPXZ79oJpg0mBdT86bccvyaeJHTEA5INnbGVAZc/WPQ
pk/8cEakSsF2N2D+N7mVFtBkk3Zh6fAkwUYnWtPuDqk5QJ3jsBCbKNecMlAR/IkWhclxwYKgQo+m
vQWKw7kwvVlOGuIHXHDUgfRi/oaznU2gfsR6Wgd9ZMLz9qsxSH8C/pcBC0BXIn5DuIm4rWWiOrCg
SeOaiCxa0xPUGYFHxdlrevFfqTB3jDqV+cDQ0BhPgEa0Mmpds17/YNWgkN1ovC3/rxpcqTOvQCeU
f7EyGLSHzGyQeojHhfwLllfgVrhrX0gftw279tFT+PR1/dIo/bccuIYfKgvxg3Cu8BpNK6Eavqm6
A7jK9OrsAnO3SbUVy+6YA+kzcb9H3TzPf579WOUZs3PhcPI7N8vwbp3DixQEZyS7O34vIrwgZnmS
M+JzDv60GQel5FSD3FvAumui+TlXsPXPetTcpB2UU9/yoVCyUlSxFrjzw9bDhymf1kOKKhacPbtw
P/YVPxso9fboaRZAjfijAWOgoUxUpFFO+6bu0NUwyv5+E9E0Y+pIX0tkSlGulrhfNtxirz+i7Rg4
op+srmKp8XjFGTPMgzKF4UhHPoBj6oQSBhVZvpPtlFWaX3nJtuimWRbGRkxqUp2aosVIzTTpzCl3
OJJ82seSoXMH4Ky/F7UWVylkiyFl/YhTwHICEkYJp9PUMLCg3Cv8+gKJ4K91TVWKFrIClQbTA9fK
ot8SM+gjnbVwJGdasVjrfAoBxEdmQalxVI6iP4duxXiE5xvvrD1JJ/wufYJ2YlY4JTRao4q/CrLo
fjN89PcXud42lnaEVFK9Gb1LDKIA1awwKYJOWc0zihIvZArRQB0oD+bIGxtijLkALYFcXKeu3PBr
Z4vwqaaTEFy/WVQGBOwU5wbR1LEjyq8HJE8aC6RtGxwEpKLR96leD8KHtywjZiAwrswuTXIKRyzB
QKfBWuowntVn0ZExNazBdpS4hOiZTQtqRq52647e2gzb5f9Yqlj2oBvpZen9ywtjKDjnRcJoumMz
cFL1S4isCbYrw0Vz3KgJcdotjTEmDMvrnQ9JanSHRoZxjup5nj7XPstthHcnhjHXToZMp2+sPbhX
GsGpkfypkYUM4tp368/o48jFeh5r7mKWwtFGi0i/u3MAo4fvVyBGfqfxjx3V8Yq6WRPt9bvpiP5A
pE40hS01k3lLMfLsaw7HyY4JtJZmPg/PMVyChR//zVYTYhp2TVcE/jJnAY2fN5M72nMpez4Nm/3A
xdkUefsmp+y8EZhN27XNKBKxUCqLdjN8My1uqKA4etmYPwTYbx66yGeMLvtQva/vYXymeRYIIbTb
6OujXFwZe2Mkc6eMovv7IZFkhUW1KOBKETXKFrk6Z6WF42YFvD2cOB6TX+HfymhP+/0P79FdgZ78
W/bD+jj1MYqMNF9uJXEnnPriDLuZfk3UxeuZ0KvnuOD5TRCec5RIuXun6oTsdg8S3Zed6BLhI6Dd
bRfkOgZcw2PFT8QsVCpUyhzIfgJsKcTNtNxW5PZD6vo8gczZ7WYrQmggaT4nqrnInc0wnhZrr4kc
RH5W1vBP9IxJx1sIB9vbxDqwuG1fbXp2spcA3L7FgYGgDfllxAXbDR4e3a2ZjzbDRcP23pgLv8Ts
cMIriZnF2P7GVgzlv7XyTMz8brnG5NdlFmgStwkCPEA9/OIEaqygbg1BJJ/ALnL+l1IgxOKu/JVV
rrylZmMFEdaDLG7HzR6tyXS15iItFE+f4ZaREkA7sFlwSWLRPDlfQQE57wafKuG9TLYmccaNoF6X
3N8+UyZzbXa1KfuAEeIH/1ZOEqjV5D6PviUz42p88k7f2S0Bjn5ZcnGTcN5YWm3km7clf7TtCva2
235IG50QnoaEN+lvIeWIh1UHgK0LrRNjLYpMG1f2p54KbWJQDDU/NRpgDtZFvBIJOVbvRfZ8VTvo
XjjCOIP0Lz2eq3bR/KmfziL7CuffFM1OhuBiayNueG9t47uZJWb31JHbbYJM4VD6OvmfgdtpDFc2
WbELY5NQitfJ4ZsJDuDJRdVIABSMz+5DkonJwIVU6LuIEdpMJeXXdsYXPUVBvMtasbjxzSn/Yl8L
Fx8kEeyrwxfm16jykR//gdrPfpUjuSld6g5lqjRMyTAXTWgJXiypiePlC8njjL+wyKvkkO0h9Z7P
qEYhHeijhHHaYpv70teSMtkm7khoyOwUFuXPDE/2m+JeRuYRA51QjjmllU/l0Z8RHEV4Q9cg9BoV
TKXbafd/Wf/92ZkIta70MWW3HsAmoEd9nXGm1E9TXmeW3Mzdh09P6biG3XHyT2ICufuCL8ujIhXx
mzGGVx+shsha37nCjtwgraQYwCDDAn7/ixMNqi8ziqGLxF7izIi7h1gz8y+QZIDgPTu4bttc7fLP
C51YHNVDvyvkDTkzbGq7nvXO01yHnKWI73teeo6e93wPRQR6/8lpKKk+D5Qzy5FiiTOWjtkNVGkL
UDu7aJ9dIwUdcXmu4kvH43Z9EWDCb9tNaVjcI1eoF3VhSgHRfKYAaB+s2mBVsJvLUTlxDfkHbnR4
jJttFk0e2iGcVm9LSVWhqkZEsEpxSD8Yv9U4rRiIKC3kZRRHJwKbLlFWluxJo2a6ToAvBhJiwmb1
srBE/swOnhnK+3wL1CmYNaVoIdLENxzRGn8uKu9qk+LotTnwigVNn9rcYodbBwDUrB4/CRcbSaa7
2J+2Ixac02253dRXHH/2Xof4/c/0T44/m816ah69si9Omo5pK2eeVn2Q1+itaNPQ3CzUb+oUObfx
vK4G9hwDxhi13d9yeT8iKMPk7cxe++y6dRDhYzEDvmrW6hQ5LYg1Jun61egdtQmsxDj8eLIHzQwx
TTgvQCU77SX5xYdLov2EKrvTvbJXdEa3sO9StGZdueVnj1uojdcnEIPcrpYhxlehs/rMgqncV1I+
9Hc5xV6onmdyahpPDk/qaETLeeX5glcRjrXtJj4HFTSooHdz1HI9xf3OkEwax8Hkkj6ytwsuaH7+
q+1wzbY+QkDcEnVlFLdy/I0FuHKEgx2/GNSIDB9gTCUGyn85084TBjFnairuU64QSpQ9nrpFQOaV
94xjkotMXEFRkrJTnEcEbHlIPIP8A7IU5w9F5y1B5nameEZ3MQhTszMLhFrDOKZVqTg9mOG3lbHe
KgaNE07RVeXnmMckyVBM1Bn5hGxzPzo/RKqSHox8tcXeSnbYXi7UK12u8fw1vEROdB3vdjl6QLxG
MIYsMySMgqHv6JmXlfc5OHI+ljAwKgNyl5SthU0ngBbv/ykwRj0QttU8HzgzlNmYSeOVlUc6GaIP
ZsnOz9P7tAOFmgpu049XRhjuf9oVlGOP8ZYU45M4bLP1HpfNPdV6Nu/Mlm+4A47tYQaeR2frONDr
FiHDJWNN6fRWq8dUAVegCXB8ij5ns04MfumD05DAmb9YnEpD+Vg/5kvruPX8xbSXph5ANnp1goWT
Hv5jFO7jCv2GRwtFhJw+WekeVUSWlhlTQ12Btw7twpfPi9hmq9+EkZG2I2G43jR/ZHuSa9+K5hV7
rE+UMCgvWZgbUQzrDkLBFbAjs+FVmaAuizTqMo/jEkzhU0KbIwg7hBW/iPcUHzZhbwspNn+Mk+3i
ceMSifwgeFt226MldUwZ8iIZFjiTbSQJ0XFcCY6oJuhdnJUICgHz0mDOVahWDmmol+K8gZBxV/gP
h6MQbO1M+E9vqkfKIhoYrmLUhll1bq04M2EiVxljzkmvryTwrV4sP9qAkO5Ni3CElZ9zaA6krOTA
xXvt+s3iEZRbtnf1OvFs0JFzIpqTIzAd6VGmwyl40c5N24wkZSl3SNT2iz00OshJe9P7gzPteDBz
OcLsYCq9KuCI14zNcb42kgyvIuDw/8egCokW5U88mGLqhS6BDqSz/oU240K3zQy+zIB/GA7Co6/f
ixzqgHJ9pszlIkpr47eXS0OzdbIkAxO5OzJt2GODPkzewMs33OzNXwMKA0wbR22+MtikS5rG9dKS
6D/bqU1iVOE0QkVX2makkWk/yTp1Wl/GaSi+GsKOWNmbAZ+VX8Xz/3xNnjqmDQW0jF0W4Tb1IZ1b
YuvoHAlPqZv9Gm5h2aUSOgiatukDQ4TcgVpm0EAIslxsNLRX2je6Wi1ZkRbcTNFXMuWZY9cggpVr
i1I6PMXD1Q+Xx/EGWlCHjoLpkDAPopPoMjq0GRr417oeAGtTjX+JSbrWUv1uJSNky6FGANl5ZoiD
KjQoEFBYnf47c1E9DHrPU7tz5ahht7vdwrHzs809Tb9eCf21w5bK0aaFAH5KN8bEKwxklGrvZ8f4
epC7iY9Mr0qQU7v0pKhQWHr0wMX6WWjFnA4/YXzu18dZdi5mgT+wxRRHJ/pOIbg6mTVocTe+VUDt
tNU55aLpaEb1RNbkBiVo4OMiFa9nSGWsNSavz7a+lGu/BhmVdRB3SAr8IB7eiEv66yiXplqmw0OA
3ZytliwpekFqX1MsxtABZqn22f7e3HcRnnlgKH14q5/VH7o92/hr+4RNprqybArHumAawDG3Cy3p
vwAsWzelUirq1CaUsolmCbLVtpSpzTY/kPpZ903m8SzTwbNNrl1ZWsQ0LckhwTQqGfVM7XZPda6M
BY9A6kRqSvJR2w9d5UMJvzWcxz0ccMZxlXkmOw6nbrXccnK5ky8z9OXibOdMCtSnEILiSiov9N/Z
awZFQEPduEtbeJOOVHA6RwUh8E3f9XUF4YnEESyO85WnzR/2poebsdQKPhej+BVEuNw0spoxPfAm
Gs2V1dp8q/Fj4rEPcRZ2D6JSuiVAh9R/Jswh6lJ4fX9oJGS8Cmm+gOAa0hJ+SNMq8f32ukPIrnRw
zxEMzhDeginh1MmJFDLQbnjr1vRO6neWb+JXiqXDqG7bnQ3NherLmP0/ylLYAggupLQi3v82lqKZ
f+AyfplEccFFtWdIZWAkiGlSGHN1Nx7Hd7bBLUv7vcfkXLVDtTsmcWS1B3dNVoRznR9jee/qqs+9
ant+E0xFVZmRNzYRbreMxb2kWvBc4/mbQ+7mNeI7XJukhB64sW+b3/sWZ1MPWrNnxo1g9ii2WZjr
0kijwcj88ZqMtctO7Yhow+llOjwTMEF+jzVlGQI24E9/1XJJ80Lpqt+9er6P0knowNeluTp48Y14
rjVZ7XsIfA9XXWdzMcLSZlpTesW8yBxfzjYDecXhSy9KVETilXxHbG9Lq2SWdMhYDcdZjVEEuZUk
hFYD07CH6eRSAfj7o/HLySvaojq6Cc1LhpvRUTsDTN9Fg90VfTfNYyao2GU1hydDIH1BkW5ZQl04
U1k57wJlcF6I6Ggq8RBv95wcwk9vVBbtLy9SvHZcr0b7zkBmz9u42dxzlc4rQ0pZbhb43m36V7sc
3M/AVJ4Uj6ZtYI0gpqGFV0cK4maLsiePc6pKsSvRZaY8RCOQ0hQc3Rs9UaXPpYVa0rqcdvxmpTNr
nxHQpsSePzrkNr0YAJrHFkgF2tm+/rJOhyqWY6GEnrpH+LGYTElFgpmHdCPzuenQ1RMm/78TZGK0
dpi8gcymbMOrnrG9/MBhcdlZf8cyQ8irp9WWLSEVxFiUjMP29Ch9YofJrGHBJiPkbR6ImWS4//Zb
CVxthN5u+YP67LCTMAWouldAU7b8/hnTXVfUT57MMGDNgsqjxc1JpjM2H8OZgYb8xKlFf4DYEHdq
QjIy4/5EObXxajiBso7h++OxIaLttygllbPsS6AnIH+7iIWpMeQBS8R0kfSSksaOrFYiCK1BSaRB
gg8YigYMIHkw43xF/BKxNPzOdTJlBqfpk34ridTFv+P2lzc/w2MrW/SEGYcOC2tE/omI+gA9ucR0
hIfD2DEL/Djica+6rAEUqLc88bKnzy9Ii96Jfyf46z5FQsjJbU/2koi+rzrN/c0ZGSHl9tDlNukc
bzLPWzgCNSjvJvK/JgWBmgq4wY4N8mXvBdniK5BpUIRmmU+jRci81COltHoA3U8+it17kBvc05Nm
iAa8LhNvv6bD7+2gvQUeAp+cGYj6JiEG1YLgzGuI48GvaJlSa/nWSonus3MrNDLUyjLsIAObhOc5
fkw2TtA68k3FRmGzMYlgpbbmeebDlPvoLfeLzQ/KbOu6/LWEAkwuIsxa+OGgdiHPfCmPFKWlfamU
16kX1DylAucZdwe0qfZfBzs38Ai3ChMb5en5J1cUQIQ4X3VCXSbcuNlB7ApVFOKeRMOD/ulfRLUU
8RaUf2T4G1OaoKz1Z8rpDWhWqSbnxnI/usXoMfcs2HcpJpnzzvni++FVR9vy+ODfj3xT6JNATsdQ
amaN6WIYBo7LKxDoGRyUVl86qv77yXvK7aUmwT1J+7kd29tNEHQsjWWF5YIXqAHvqYvIxeIwbFq5
1IggCRHnNUbRRnz0C/3HV9y6iA+Xnt9fDX1G0PFpAU7s1DtXp/gfQqEZ1IokFdQW1h/C5Xu+29u+
bqLq1sJYMcvl+Z1lib4qbJTZNWN8FwD4bL5Wy+hdFMCyzxMduldfIDDAI0+VkkbDcQbH9501k8r3
Tji48WU6TSZIWXHWx9Eu7sfF4M+GLotvoyX3tNxPLDjYgth9HAKxefy0LBna3/AYfKycyEsSgw4Z
VUypAUIhm9jXWJlQIx512OypW2xE3lg639/WmlrljkN3Gi7fKcXC+KHbqsFWN9ebpUwapphMF3e+
VvEtrdX1jXq6jZiJixoiPkMccKdgjB+3sloEQs5n5C6ay+djuX+EmlVX0KveFT/4BPjxRzWGFH9G
hoeAtoLcnNi+TWupuG0BVPcvSYqdRFwGD3FQ3QpMWd6AQFd4vICnKcvAgLhQIZxazPFewAId/CAF
hyA3yhvmo3nW7LNezbl8NsAhcT9P1onHoIIO3kbZIbssxMtHpgH23xxgulCfjas7KpWu9WpDAzg5
vqz27B/9JQ5c8u5EHj4U6ppKUBZjzJs1JccLkOkq7pkTpG6Baxyg5sGMhuwdjLPWZudT9B13/56/
4/yJhiIIhgLhhRDWjUpBtZWi/DdWIcHopmh+Z5YxAh+ZgfU6gvHM9gTnDikAuFU2oOrMc7bE35pt
utMy6IlRnrJJIlzQEH6zJ5//EJ9VBp+KfbVozBFhZGgykgezHroYYXoJbpngtT2uxQx/09Eq83QT
YqwA7UNfXnaVuwTHNSj+7uDmFtehid6ZARv8r+gKhKxoxOKhJVJy5tOl5dl9QEVtn3kA+b571SgW
hoNFE5GAW3kJQfLthi1LYVnndoNtXEecdByRNZSfxU8HFOlj/l16n/QB98mxd2TzTnXAz81oxbtC
KwQWsp7UrZXjWUzDiNpUijYHiLZoZQf7N8KVp9/VFf+6uU6lWUKqF7lRIWv0dlPhZLYU04cucJUW
y4TA+25unkPzfBzwYZ5GXMjcQkTwuKNihmgwDOZAgsczwNDJ3oPY8BzzihQvGZql8w9wT/6Qm4UZ
oaEnQqA/6dWsU6/7ysn7VhwRFXeGS5vRCfhU2jT9Yrmc8gXMbw6jbL4DFDpUFm8sLcxAuzVycWpM
ACTUJzvIFnOg4P7fm+tgXtJlCw07WrXBJehT07VHKIMRQXFz0xrCFj3b/BRt1ozed/R5nqSIWcE+
UDlZGo6U3SOayxRNKqzxM5V9T3H+ZVMUmizSISPZtnZqIAOnH/wFSabRJTPldIkjmzmQFjnh5mKb
ujhsBq5wap0QRF/TzliIqsGsCJy8bMbK380FbqdKW+8KBJ91qrAqWI1yJh/kagbfRnpp2EHiBbTu
8DAUuMeKmfWpTjZM2YAF65m5RxAHII77pbBy+KFCBeVDbYVXNemPIc643szGCXQYLnbpzUjc+1eq
ZYvQ+2c1/MDRwOKKZsscC5JMQbR2/Xk8AHJ8d1Gh0zvPdqZnGrEwjaL+gRnRKUusVQlsvlNn+N16
M73tgnYOIXVQVPD4k2xtOFhYhnCrcfB2Wpmyvd3YR5oeGMw5UJFctaNkz1pv9PTkhyxS0f4l/pyG
8H2p90TavYh6v9e4ZvM4SFkAIuzSzdRW/XIFHKW6EMUg9Ch8cQNj+1H5IyWmeI1XjcGL/xH896t2
7b+X2588E/FbkkSExJ2mPAVSW5GHIA0FRE/XRwY2OOnd5g/DUcpMuRSrJGCMNPiYZWihRccMG4fx
i5v3Bid/KpmDqM8d8YyYU/6cialRHfP9L670spmQl6qZbTv5gJ+E2yYp7wKBUd1ceeTKUPa/atLH
C3BULTrujgdq3/DZFWoUNpF7ErQfrztKI4p2r3NsW/mhgceg5vswKdAf/gR0VilGaQNXD/ksB5HR
cn0P8KjuCbCJFQHCf4fZuls2fJMAqQFWcxtv/CfReaUaxQGi7sUHV+fTFgCgjpQHQWv6mMDKBEnx
MZi6gwrBJIVYDAMdniqnWrxdN2kX8L+h3H5d4/Ojoj5wCz+Up6oD015oRPIwgKtE9KeNaryjd5JD
vX+EoaL7gJk+1SHDFuAD6oYTtxJQhrk57xE2C3wwMdiqasmI96U6zcjSr1jD+juhysShdTa/zC8K
ttBsT+S2ZllJqSveYSTy2L7AaecxGwmNXJ9kTvM0PXJk69aBluvTQ2TiEgf/Z3Z6c2ltKhAWsv8K
QOKiYm1Q4ztxvBuRNmXzxlA7kH9ulsApJ2A/cWh6Kh6I3qPnbwo/NApVIJdrn2rnXU0Qz0efiVb+
dHi/DzZp1oq5uQjso09iTc08eDIxJZs/S7LNv68+IsKmTD8pAXDjo1eId5twjnMxK9pdN17h0BjR
LJslkre6Kgk2OXJcKW8/hHLwMY1CqMHNDWEucGiRaDJqA4WcStGI/i5W1kYd1vm4+tqIMzgJaF2U
sTLJV9bUV732GUQy+/FaqpOK8EvNOW9W9vZ+xLa9KgnqGEOnflNne1YwRYNmN14M+sEZL4R3fgQi
b3qVEMIcfxWhAzNaF2PlYOyB0Xf/kDedI8+M08HgVaCK/PBgpgvPd8hQ30IQtznWHrI4Ziw40/GJ
ja5wL91LIdwpzo8vyvpc+o/6qq+QLtLoeMSljtxmGwBssH/+mbTmnNAvcq6CM0QmNZRhRTPM4+v6
ftD+Zy0ta3pP0YqV6YW0oFtn/79k9Cb4JNxyr4gQDbGQy6vlFDYV0BrjzFZj+q54nEOgSzUNWdFv
1mHJehLX6pBpl+t1WIUwVc20SRnRg4DNZsEvDrXM2DScSXeVEpp1mYrTpGUUsR1r5Xz087qzrxMH
cX8z++OpYf3DhzAnKddoOnPKJ3SiIksnf6apweYxmpSDEhPsGEdjILgT0OCSXCANoRtd7eqnOXB8
XS6ib2zcr0x4yY5Dpt0OQp/nBYcEUmCfIvy/Ho7+MAjNLaoP/G4y+l0v6kokDMorFozn/aoW3k6U
DxiIr5b7WecqdzM5fteIJij/CyDlTq/TPv7KqdkAgYOpuyV28EZXINDwfQN+H118+yK9gpFCDIzd
HOGzRS/ERcl1DVAXg0gf4ApZa6gAAESaKl7SZTjlXQUJtSGNcRxZQe9m95e22mXjGQ/VV/Q5C4Fs
SByMPBF6qE4c6YguHZJTFcSYIFhiW4kixlf8aTla3eiBeLa/eyed0ojquN4mWV8ksLvTbFg9No6o
dgbciNWtpOtI7zEpf8iOKHmnmmcUMza7xYfSd3udePt8XYIVFDBuK43vDs/Hk7TclJ3ZiOm+i/Zj
uZo+dsnh9Xr5lbU1ljmDwRYrEA7zFcBaM+8H+bmuUu75pqlRgwvd7No49iHtQvZBao8VH9bhyvfa
XMvSpUJqb6rGLw6XpPz4w0M+bJ94D0a8lb0zvcQFP70A2UUYWP1BHNDFILZTUjZ4BPcRSaxQWWPL
glH8aX9veNTFYscTuKkkQycQkGNYdSAy2a+KmkrLcwwQJl4O/rMXywkdLd13L/bl8Dm+3gcxMzQK
3L9Dj+R00hrxdGEKJG9wFpMXQcDS4Q382TU4rlHuMWByJ6DZLN83LFnVS2X9OGmnjwS/XZSgyaKM
b8ZqhcVf1KeOhDP3hUGvzqg30Q13SPCl87I8e1Ww7DSc+7H4NgZA/Iu7eqlKsLMjlQtefxwkqZr0
rfgc02jPBWpxT3EDYUPR9ocjtKZwxxUWAe2XCraI4rj/vTixtuK6tpFZN4Lx7+tDv+zq7pJz8w3y
yijK+3PkQGCts7ZmYTtTHS9T1EmImZIQ/m6JGtFWS4Gbeq1mXBZaVL0fsB3uEl4Dhj8vGL1YuiHt
NCdKqltE5cmo6GK/1QSoIFDKAiXpO84U0XzVZVQlNu+ZJsHFtbltN6QFB3JnHcFEVmCyezUyRRIh
nmxd62d1I1/OcsOIuGWcXoCHYMWysrhcGfR1bC9tdkAc344ArKLc/yJwaDn3fvPOFpIqTzlaCg4/
ULvMdUTbOa/k18xUnoV2acGPb80BHG+8kwbQWbV9W/PcZjgmBAS5Drbdrrz9H5VSuX+6Vs8vMXqq
KvwsFWtT7P33eMCpBmw1jBVZDL4UHKMhTgJbclPh56gpv/oGZYdaQqOYu1FNnPO3myrWqM8h3tZ8
zipsul/gLc7SMPgsRuAIsPJA48OvIeslU8kjBc05+jhiqgndgqN80bPyMO7lJheHVxCf0z1imUhL
Tz+j/wSgbikUacMiBya27fuI0EaJHJ+zMVQJQJvOn8Vzbsdxza/LtZgh7oMEbocOGKMG01uf0jyg
FHhkx+TpF+yiy7YFdO64AtFbAM70HSW/GonCmUxe9zWzXiUD85o3oXlayx2udDIPauSbfq5zvnoG
BEulMQRh00lhVFtkSp1+K5ddhrNUaHJuyThlfJOtuVARSKdEXt19abwWTAwNI98czKb4o6w9NNIa
4wFvniat8jVE18HOO0/eotGX4TXfY3dOP2aVzzEL59szw1DoA0CB3Rg2Xdf1ZN9O8O1BUUUI18JO
i0/97MUmADIXFLPAb5Ui5K3QFWKcgSn1OLleHg3fIeSmgrc//jK5ZupUhKgnKSVLFPFAId0b8qyw
NWyPUo2wI1GCwK6k+NvnpQRqtaRcJYMnp95zLDLdK57Rsri+l3lTbNg3r5HO/b/mEzSWzLfkijXd
ySKMqpKkUFi1sfNZNs3/Iu2hoV5M8O0QgJQRdnXaytdQOdemc3vmU7dXJXSFOV4Q4emppUceqq64
fJ281JiHpxqiQU0pSoT5hH0t2OhsxafgyoNiuceApaAvPlxz/ueOB5O/JynKNDn+qedFsgKZfdgE
FdF0cTs5WLSTQ3OzvscFNLgGqVjk4m5le6Ot6wcOzxN1R3U3YPou7Aqo47U6n51BWfBOyMwCq+wW
TNhuPDnSjzpl394vegG7+jswxcfgY8lAJ7IVCtKUcKqfGaruDmLDlkbijP5SXx6Cb6uy1V7zzLxL
ji7r648JKTbjzC2sZG83Q5+l3JHP3Is1OMQqEjWIZFGQRtSbxvsF2XoUFU4vXkuxnsERWy+XKhYs
smtOrodvtsvdSKP/szmTSQ1hxUOWogRBaqwlpEU91o4DqVEyQjaT3z/WnBWTLcrDvNNyYC3ssAu3
onBxWmbn+q63khEUEO5xozeO9o7EKszjR3wc/Yo1S6T18uv5EW8Ncxh4tBP9pkpFShH2Fq6UMvLw
S93hstQr7V1PtacCDneNLiZyZBIcHrWm7Xeo6C6nPcePh67wcnEYW/65VmqZ4CyZIGjMcWAHRrAu
T7zJN63HwvNONY4l0jZIVdupIJQLxg+Y9gYXAB4tz9l/1awhL4LiTqAk86Abny2ijw+259z7AZfS
VXUY3uovGMPMrNM5EhJyKy1SMNO+oRhif/zFoUcnH8p/m11HmGdmRsfJ7+mmAKnuAGz2nQrpB4it
JuYcJY1AbT+NLsUsqrQ3jrjOxl+Ao+U30aJRloN4jPSexLX/CyAk52CerxJ4WxWWyTRk9Xl73tAH
RptLwMyFT2kHZ2PY9/bG2wszhLO/EF4evpGjFmM4nHzuaDYG9hPophVZcc97R9xpTe/2ik493vWE
oP2pXdNfLPv4BKLAgnqM5zrm0/XhBdhww4q51YMoTMs0BcvpGM9vvjf19HIxEDZcTNWVaTeia6OE
HAgeVUP8PrKVIQS9YwP1UU6ye5ZS7NcU0kIbDCsm2Yah9/ts8/Ri2ok6JbkCBT2ThgY/XJmh7hlY
+rbV3HifdyQzpy47vd2acudx/I33VG0vqIWwYg12o5FrrJB+o9byv9e/GlbqQNwCRrhk5UC1i0L7
1puOzrYWjZ+bqGpyJuQKkwWBPLV4KO6hVp3OzufD+9SvkbpOhhWLdbXcd9Wzlhb0rbPXYU72U/F0
Vxi+pHeAPAKjXi2jRNze4vzCy46Nvxrf0pNhWBSrxI0o5+9uyqxoAa7NylHCBl9Lh94+8z5xCHW3
VnIPb4MLmjnAjGhFX8cBcwRKuQ8YFOqAOngfCEmUgTWccfOZKKMNMQKMoedxvJntf+PV0iJh0Crx
0aXrU41FRFoQBAabxPNYydIUlM9bSURWMkzSNmrWLc9jUmjhD0C0lZyfwXs2xmyUa1I5v3CvB0ky
3lX/6vq/g+gqCZWiLMCu4cQhKwmZ6WHwxwBRDWAEFtMqt5H39rwVPJFzhYV+4MvYIvMGV0ZV8Fpf
HgaM237w1NyhEK0bkYwq7JghFFirbmSOmrMiRQuT3iw9DnPPoCKtYe23fIrAMpVcSw4cPUd/iMeI
Q/6iIzWvte9Lfx41ZGl2VL/KIGiKFnJMdHCtlFhISubnFGmk7N80zQh1yjluf9Yuq9jQRpOI9wH3
ya/8kp/di3LlP+Xa3fGHTMBDd+wFJUg28AkvZwkZ8IqB1s4gOLdR1q5sk1s0QyD1j8NzBy5AFm5z
lnGjVMI5GtC5gOcZQw3Ot7qHJFv/bDBmfR5n9Zb6YeoD4NFP6BW8XVoauOEBd4mf+3nJeRi/vjFL
Ogs1QfnD1sOkbGcyIwXxUtk/XVEjBm+j6hUHWCQG8+p0GmJx7NfndqmFb5ldEiUKjTG5e0umg6ob
zlJGtvevd4FjT4IWDRLfTpRkhvVHRDX/1Wv0m7pFd5mhLQboATZOq1VjaLGf959QCcmm+xugM2mE
YNjhB5mGmT7DCdzktyRf0Rq6wI47/rQLOIzHYkW+xvKiNBpg3sIu2JEwqIdIOdHtlos1qVr6PN4V
R3ourb+M/krRPleIBNdu5RUDxBfRcQ38EWhy4oAEAJfcXoKE4WoBQiYMkEvvDkWsljwWQTMWfnqN
5gQKHNvTk9IT0djjHbNsggESP236YW4UXY2ykSL0FIkiJj7YI0KAUtDXbaKQG7R7LJ35KG9qwlwu
YA2u/6tc1YK8iNiSBONVtwG67ENY5Zz4QLwrHlfDoPhxTqrIslNtQvFFL1xD7CsLTsE4HPvdy6M8
olQL/QapNGcvjhRwgcdG+raupgVWzcAzpN6ezA/8btrSBmXk7V95MGNzhrQ4Mv5IS+FZj49OnVgt
DgRzifjP6gXJRHCJoFU0JPHnkyns6FJv+h0WLocKyk+cqUMztDbrhJ5he54DIr3euy4/jAFsSYN5
m0vCY21TneZW2ZDzjo8sjJmDEsb9SGbyK1pYzKxiy1DirVpybzYylMd+nuR1ggu51krPzESej0YO
tFS+qtRSQzKZ1z15t8vSJtP7u/+R6jlYIXIrm/1h089fIDnYzEvcNrHZchlwrIEISX3ZFias+0ZQ
Oa9BgXS77T3ZKl5m95147UsF4J1iScEtePk1s4li5vt7o2chZAaZjeMFhNV9IR++H9BcjwbSewC8
GCKHiBieLaxyeDel0xnIL3VMsD4OdLpG2qYCEgOmr0ONrAQAF47Sv/W7OvDi+ov5UGnnP8Wnm3aE
nMRr4oFx6sFLfrsidsofsZtA07qM9YQkyyJCmAxiTOsiT7gTAugoFnjwoO1tHeQ4jvHv1/xYt5f7
cmYR5B04Px4Ey7zieD21PAjmvQLm6hl2rd/F2OXt5Rw8cPvvd1aJd+6bSMgMh87QP5fRvspreAm0
PDxtRPphLnXbOkPbgQPC99nHhBqsHLkHGCdFbTff3w0y1uRe7QwKv/mQZK0SKgIcrGQC7ErAmOmx
ft4zphpsAY/C8XbC08vMqF0HLsGQrhZjgYWUkytZA9BMb/j0lQ82QTNekPxNiD687pDq1X2xtbLF
lHzSYdlVkafKmo0qRcGbdvNhm5ubveswTI5nBmhAtNGimPB9ZkGbQXR35NSRW6EV89hE9n7MGyGi
6nDslpbvrIxzsAr9ptUUf3dFiOrZ9PwPZq9HOd+9rKwFaS4YG8h61KDQDkgHALTWN+J5MhAql7wW
Y3CQsT85K7aq1koloB0xT1unbn/qNcl6B+TIxDdTYbIdU0IMiYv5H7EJxB+537wj2d50a2EspSoM
sO4WOKIEroetBOlGRb+Nw1xhTJESoSLM9jbyKmC55JS5TeIhLf4UCwzFfIupO4ujb4ybvyv4VImp
ZMxAaWkUcUmhbg5awrqcSj8mxDQYRxKvQrt+Gm9a+WB8oRIwbjuyUZQnkgc4+42BbWoIC0qEeLmo
VwsTNyZcOk6cCcw6dQ8mq38OuPF1noNu4p6Sdxz4rOTsywunKUFXYToHPHI7IZBWCjJWxr3mrCz9
aQmYcX+5wjEiO4j2heCnRIXyD8lQXZmDo7mtJCalQBZp7w6x17npPcwg38WFgdCtxVmPADSid3R/
mUGMlwoL6iCxQYkOX1pLo4Xn96WUTyNDWbK1RGFnKBe07YnewF/V+uEne4MuqIDtDkCMts8tSok7
IKebVgoIIy7nsb7zXw49D89IpKjiDxMdRL4JvBHErSYLi5FNnD/4/4pzJtayfSE01ETLC8e1/nG4
NM8ptV+Y7pel9QaltjNfTPO2/lV8fuydlWugtxqR1QuIKx0WT9EIgNIAZvjHeBrnPkmZKHQg81SL
qFL8+SKwm2K0SMXx4FlXMopc99dVe1g/g1Rmenp+9Zu0dHhDWyedjQjWFOTNzK05Ckxi45THILhl
pXbC12y4UAeeqolq0K1if8Ac3wu1umlwj+n73xP6wl3aKdaGt1wOs5E5z8uyigcTFtNhHiwYsW2W
TGrJAnDq1UrrKfcpOT2K6XYsT4CWGC6+Ub69AmvmtwzHJ7ZAZSo14XDVZch+0DIpMBPqKhNVL8c5
Z6HDCwAgBpT0k2oAY8SEHAXgEZGrL1WKrHvtTwoE6cBA7IRQY06UOo4iG0GbEC+0hgUdh5RfIl7C
6Zkvcf65aJcT2KGXUTZpPJCac18XLTFCTDUIOdPaidvFLY0CetqGEjh7LxhmHtsduDEI/BTcetiW
TxXRP8PrCsKZEmD+APeaY4CxxoWWn++paZi3T6dKQMuzceu+lrOHMSI+WPYNBOXi9+zNy8KQo7bn
5AawsP41Hte3V/4RJGT+l3s+FmXIEVKSbOBw8TIJvsAtxbIr3+4/q3G3kXETikU2ZIFWfGW25jWu
fgFj24fRVkGxACykCvQlTwNn+UTIJQMTZV5QR2P1n2V5S5FNIO6ksX5CoNj8P+TIk1ctve3lI3k2
fpr2eUiKXSRkgebEoG09XeKP2akdOiSqXuoAixDxZfjVFUqD2ot+Os6duYB1sxJok8L+khZgiLhM
eEUbM6nRK7KsoD7LbY8IGy1P7gBhdMxR94v2yD7kUpQmuI3D3rIhqDQuZl4BJ8q1bWdGn/c6MJXh
IXXxobN/tGPUgKAHAJ6V6xACxahgf+yfGOrf77tXsH50K0BOBoySTL+wR5k9C4C8mz2HSxH5WntO
u8dGs0YiUhWvrVJCHxbnsvJcLKaeDz3JF+wD8l/5F3lzUTWUKkJHAGpFQ1GQa6Dakj4Zy7LkDCpq
I+8nAcVZVUDnTlqWp9TSzmmW5H4V4TQXC5ZfAztkzRZsGt0+hLTbzoBsv1Q4wwK2jZRiNGOm3gAN
/jZTu6ur/+I06DZUTFcmOP1vZtmUiJrbrAbvTGGNogqdiEUeI8re902XBY4tWMfcQibKqFXV8gd4
EJgojwVxZKZvRJIPLsfHL4WLnYc2OH1MbTCLkGQBw0MPHPCp5R3wg691o0xhZ1cbXuWp28mKldEC
6SRbRLK8QUd24Ubg7V8MGzXB9a8kxEuGPObVATlrvGqHNnurFO4p2BXpgRUsxmAlU6ltKr0za8OU
JO9QByJmk5IqbDCz+rdQxfKCF23h4mZ2jrGtVtHCMABZui6O/B6HoUTyZg/uCkV2NEfILQr9vxfC
3VzVEDrFenIrXRq1BIHpw2KZimaXaH/DKoR0mHUhXAYKvPqZRhnVkBVj3DjBsbkyjj16LUD/PoQ4
6ZPiOI5qX2NO7Qef6RCjkH+6ktpmAzXkxj+iDBT/W9Dekgn04xd2kgFGc4Q3rVw36gAQajriTT7Y
j22F9chtLlc1bT8Jv8axGjf9FvMIhYcvkY8pZy/xgDobfecr5xKk7kNGZHiNWYWWad4lZ9SOO4Rr
WgOVUL8LDoZOcSqFueN1pdt7FF0ZGQQyGS7X+M2s4Fu57JHC//wzW3mqspZXCOUiuHGkbnGdq16A
oi8CSRbFZRpx7DpmZLpRkJB2vJU4SB6riAEB7SNTeDTZSTkclMuzuSzAbwIEagBtAud5T/7rv5Ex
8Yiew8y+is9k29Ch2k/s+ryV4k+UnoDOhPsi9uLMY/HaSafNfcKZT456EbGu5uOMyiHn9S4zoNSB
ergrWxy16jlfxFaqZlTpLAflG8ieds0x6Ol05RO5Z1C3ykhqIbo1yGVyDtm5yBxk7AqBJHZS4Qhm
KrT/eXxti3aIKPlzWrbsXa1ozh+DfTtjUaZizEbGLwnfTsE0IbysAWMcskfQsm9ASduL8YDS+aFx
AYVJThAsW0mPR9bIo3VVcAC56VvO2fG0c3mw9P0g3itjvm+S9yWoEqj5EwAtMe7NvUJiAPFINCuz
mVu47pIajw5rKMXOoXVeCZVh08NZSi/DcvFeNbXlVzzkXfyVDwTKrjpZFJxHlJPL6dr47UiZBrBU
qYDxjxgqMOZqpq+7+nvY+RtM1cmi1rFgAlANeL7VFbAZ6Xq6YcnHv18zoTvEtg8vfL5ZNoJ7qyb0
f9R5RNjAcdl/3KcnSHF7GHRzC4aeB9XX7audYDSkMjhefHTfL2zoeBTxbKRVi02Trg0PBsThJE4R
Ht4pu+6tob/JnscWt/9xr3v5aTlYiGarOKbHZAHgmVYRowNlPTjqjVlLjm4jYUsIb1QlQkdqTr5L
TV58GGBJ/Lwy6REAkI4LHvDVWnS9QT/sFhS8TsqdYCuzHhAyET+p0YhNURJLiP03bRUs+q9CvaXP
Yhf4FQ5ZwoBS5GTgrnVO0AGC5dYLiAM11xtoabxvlS810EJyY6KGowoaAJAp7qeZ7ZNVVN+XrhDT
UO3ekzOwIm1KXgtdaJR4NNaB6uj5Ru3a36FI1iGdlfDLX6OOhLRGi1O/wZNNtdqjB6lI+h7+Nlyt
zvAuJfgob36sWcFccHPzhUMqz2nyRRJ1ZscOKL7N4jUvoUtNJ9t9mHh6J2HP/SG7TqEkH9L64KHj
5CADddoCyyLQUfvlHHHtMON4kkRssLXIn2n0nZzsW6xJGPsTicp7MfV3CNxbeOVbyuY/7yjPAfnS
IZus2VCeJeEDPNpX6855OUgF9ocEKeUqEOGI4hGEnrND9kr14Eyu567KPWnhW5ItH4zH5IdXLbpl
/1hWSfvjlM1yX3H6Y1o8YimTLmU1nLpjrf3i4Hx8XrBMNgYyHfL0NUx7dmDsHKnrqNFZ09KW5lEh
blRwFlHFWiSPvhpHJgbCmlwEPqPGrWyLRpZyJXBpIQ9/E1myNN1urUJKXEwe5BI0E86bL469HGNW
W0i4a+4BCQJ9m31nXEoqkbvxKnzwyy8a9unMFVbe4HRJdy3KiL9bZSkqKfy0kkJYgChGEQpgCAma
fo/hgnC5Kzrl/nNoppSYtMBvG+Ik0CI7KrVoPPMFoHZUPXEYSnB9Rg4dHDkQ0X87M8w0ZCiLwwU0
7KVcGwQhajXmZQ82LdpZZl88Jw/f1uzDHXnPiB/V3OuFIj2bVenxlUSvwxmX5asMoVWnVPiqQ6VO
rMji/ewtnQDIpyzlRE+cEhOFXMHgMPOa4b1v7oexgKVkmbbwyyuyWuEEjD1hWOkuSOuA/tbG25Uh
93DtFFYEvWNwbiLQGwnSxOJGner2PF/FALF2BsXK9KnZSumAKcf06SQPo3o7MVGPNfkwYfnTYuzS
unCabU9Rb34FFRiLNjiXnazi6kJN3cHl0vDRp1+gMSg5E3HTdkIqi8S8vzXMfMRfLHV9fct5sKK/
8dh+qqAxPGVNPF/o8kgpOVoZes03iF7WJdrWkit1eJ2iU2Mv91ip49tl1Nc6ZLTgig+kf2hkx0+8
wQJyPakeURH1ONroJ8/drpM8fy/7boZaSjm5N63C8TmgGYDoTE5stJONvxQoj+FI50MR9ClKxavG
egh2qlhYkHEUqZISQuz48u9tUWc2rhCfOr/asPltfkWwQYhyGFqJVZlzE79uwmHJ8E7hvCARHOKp
sZDLaEqBTH57zJlXtM+c8MjvGCw28TgODR/BlxB8uPuVB7P5LcJTUKmsjwCG01InSVFhjPYNWkZl
oJm2o9hWDzMa3jO5LXDHaA+UnDLy+lEGcBupARPIeLiGr/s/4Ok/F+YZCfbtmRaE8mqBnK2Xak7J
Ot1ovZWcU7Q1w75lE7cSJNmJvzTlek/lknwawqoLltboS2lXN06VXSausoulVLTgNn2sDPE3FGaC
gaE9uD4JkZgv4gr+6E38bKV9iFK1XuwH7C+aoKtYI8sDuY6FGYPsJfiejBjMoMudQyNkUxCQ9Pq4
s5VMPJS3mtFTq/5BNaetBzQXxqLR/lixLNuc1bDkYC2bgOfrMQhElQ3yhDVoauyR60nfKv1Tk16r
+w/TfbCbscAETffimHN98tmQc+YaMT0f3B/qYjdnrbw9faQTU8xuQ6yPh9SKHVSvMTievxqShGXM
T28USRRfycXV/GCe9rIQeJKMwI3t+8UpIs0uRFZa1vo4XH4GNHZj/8BpHkdDA6Ud08Xtqskq0Siw
7U2lnT1qhgRzaf1V62sjUi3R1YQAwcbwXWmYbetGNQt2X1o18J8dawHvaV+YeoUC2GnTvlY+HVSY
uAetpV1EtyWGbOXn6ZxzsjxeeQOigu80NmPQOLE6p0d+wesQmA86U0J16ZNzgcZUI0kdYpOjaUAj
15nTfqPoMJgpkcHQpxLvFg3T87EZLVYhpVjF7Lpu/2tqi4hKfskcz1RF4gHQ2ND6TwbbF74Exfjk
fh6L5Atw/oEgzGQ8lPZ1tRnkRBFgYherFAY04FSmMFUOe42LerVIDWZpdNqzRCf+WkeycaostqYs
/OZMdFyOOYwd7KYOiFyE00tvAIB3fgA3QLYqjxE7wZTDazqtIHg9luB8cRYymTuVbeJ/bYfwJ9EO
UEHxWtC++AgMpwRfltglE0aih5bQQn5S3mpvy9ug/0628b9cIQ3gsmihkFRfM51t3ss8WGSCSTYQ
mzTyKJ1VQyxI50j3NZq4BIzftO5+vjyPQXTA6oodXIbjdgitOScw628eGJo1/Qz2zZ2CFTBSS9YI
f5u5qL3yKlQkQ49VfVb/YcTaq+mJTTl2SVVo10YpWXbbLvOJE4/teKZd39Ir54q3DfRn95KiABoF
vU5YyvL7begJWo3APjyHNEAf9W1uDIeBSeA3L0r2xTohF7hX1pJ1lOkYhowo/JrLDQ4SFiXybJSf
JQkDJP2Goh1kNZObCjLD0spCyxazEOiHZfzh9Ovi+3mZSfXQ4HIrRZCoaIHUX1oolaLtk0otQtI1
blrVdssVSCuho/EmnuH9ExKQjwDlwi3E1bpPr86JNzWjQx8pMMPkg1i4TomMTsWkNhbJC834M724
pRq+nlc+gXNJ0pKUt2M2moqpbTqCsUnM2F2oZFCVdTNZ2VCw/6FpVO2i7m6ttq4WtHQI5jpU05Rf
eIdsXEhLph5xHeqZXdeRbJWBPCObSku7dH75goOYb7Dl9E6MaBFOxJ5TcxEkCv1mBAM3nswkaBIe
IG/VXfO/kHu5YX2CFXURjJTtxfP0JTg4q3SmturT5UIm+8i5k+8XdfUHo4wADjARgPFHLawXN1Iv
1he/ZM04ISwMz2mpee0czg1nQdy/r+N4OJlHbJ/f6kZMqC6cFu1tNdYFtNCp6V0O9Sz6svkF2qHD
pavIKMvD6sT+iAboWLNrJp4i0SdRQjprcYWNNyPJzi7G1pd8EKlOitReu0fX9A/zpFYKIqCFXIdk
MLb7zd29AfxYi/2kuLpZMueEVQPdSUqbtwzuC/b6DH974AdvgN8ocaeKHBnre5Z8U6GmyujtjfTs
Xv61wFwjYTVnCb6hDgDsKvPFU/eydrSeWy6xLlLr5NDX1W8wxU/fHFfHemFyYwNZvAPWIB6/KdGV
CuAQ2J4amAcW5BY6m2XiKqTPtbTSgVruA4EcjHObNG+hIp5DF/l7fSCKIsDlDKSLD8gsDkpUZMOp
8FatB0e4l4Y7R0OOK2PaP9eG7CbJv/ZllxKQCrrysB/ISnF8WEM9xlA/llGBsS+jOGO06xoJmbPx
fsfxZpv4DYPiy7Dg0axOrZLhv0t4FMJezKNtm+Xeqy6NbASMN2d82KicM+cNxOz9Fbzd1lXV9xEY
WFSXiyczZmLzSEZ3YKLUD6gGHOB0Kqkke0bMUUreT+RtElyXjpcpEUpOqPx2GZSDc/SurDV1yP/q
FWYXPKfRrlCEcC4MFCk34065eSvkDi+nWY8v204hvOCpbEAzFef+HbHc32mBr10rjQgZ45Py13GD
peXBXle30Nfx1t1UkD/Rhd7o13bPuVU8DhwouQV5Hg2akqJ6OQDySGZ6DehtbRq83KNwKgmrjHRV
mDrfRRlM8o4Xt+63sdFJJg5t2s33+nXpr4Qtlioe2sUY2hYsc1gMVNg0OggIh/y+GA9xUsc1Iz6R
tfLzEL8uMRn04BlVcMLlgu2l65bD52AUuvMLYUhxtmOV4z/WN9wR87PvuqdFb3ZOmWe0zWSsAd6p
065xFKnvj5pQhcQIQXjDCgXyveHxGWnPg/1RXNkSY2v1ZXWy6NNd/Esdh277WAF7nXG3zrmAgcYA
SgJ73rkXexusc45BiJLUO3TVHalKnEK9ZvIsA5O8dMo3f9MvSttj3x+nV2jyOLUgz49/g859w1GA
pI7wNs6j76+lnLdMZR0ER/rYCZii6tMAdi3zhKGkHolaKLsAw64rmqgEOy1GZubnqN80ywroEmZu
k3u/iVw8lHK5YQYWgPFRRum7JkpH/CI/9qmdXOunK6B/Tykr3XFXspd7H4RSEGMRy74ratsHbMoa
h8IJdxCcMvSLqnZruE+A+5uecG5Xr6XL7BThc61NMjxl4Axfz/M7X4D5iROFqUT6/yKFr+hCK3UW
M0MRiPaeVnVPaV7es5Zj3eJtQeQOr/HNn4U0br19nifE3GlDccJiwV2PiGR9W2hw6PoZWEXTtPhU
aotl6T/ClInmMKWcMQdoHSU7J1ea+04A36hEEnmjr9hzTRKFcDyATYSASuUxBOO6/jEc8pfAw9b5
4bRcSNUg770/3ksnx5Z0TvJeXm9/UT7E9GndNzEfzlfFqe7+O1p4MDWOLtpc54rAofAAVD23W8pG
j6BDWUkP1BH4qGQ3EUskdjGRN2Nw3LNjR3q8F5nVuhOZ9QSK9fxnNnbhQZbVd6HrgyVCf80NO8/v
MpSryH2XBhuqJsquBdLbW2JkxJOlvhcICIEIzPk2E9Z0T5MV66cY14rPY3zqc/6LOinxJR6SgWN3
HAs7+kgxTMm6YvocjX9a5OHU/2V0rJDAhQshYcXgsOELIGlqhmaFRPPyMVhTbxtvX6nbvjHwd9GB
y65WzBEME2BdDzFfCGjQvoJHqOLFwepYcslM0Dvg/HG2g7kOnHeJU2/HS1FqKW04NoBDaw0vPgS6
/bQG9Wj4r9WpuBptDWo9hFlWpQEoCZC+ws7IaKuuWeJwN6hsqXvjGj+hj1qpa5ZAdVkltclijY0b
ZqEoab8FYsh5mAHKqIbWP5XmGNhT0+QnPPO/WR5Rmhx8r0jSRbREjKiixHYjVxf5gV2DyPhX8gBU
/fkbBTi+W/dEc6hrU9Io6dHwCGJjGkb5wnrD6p5eWL7VKKJLxO+N5IFyviWQ/Q5CDfwVkwDrc9Qa
jKU8T1qSXlGSYvv+kVORotdnH+QPr2r4agChjn9kRJVX+b3K7E46pfZVQP3pM3g2U36bhSlX+916
WOCAk0qkg08VcP5QTcOmWY1ZEDqY0L2dTvJWJHrduTBBOGU3SXBvT+CvYrHphZuswUl+D6b8MY7k
CU9dliOI4wP77hez7/Jt3FRqkNznep2stDuY0eQsf0WSrTtvj9pcnwXeONJtMnfE+O+0dM1niwB8
G2jAAZuMMhIQnqN7AsxvUrdtst7XjzIBNYKFp2VU4Aj8tdFgL60GHebcEWgu3lVqEBKk5JYiSl2x
/SD9KKDzMGluv62v6bUEEMWCUl01fIxZib/xvkOdCWOSaPgqC9qnCpkAAET86UFbGqWrwk9I5Ip0
/53s/wDwVZR0MN3eRnGE6xHJEkVTbwlnU5omoLgoPNUvfwfZYZUu/00fbpM0JidoOyLkf5xAZpR7
j0IP6EokIQYkApzm3TcjfiRcOBv9KlKl/C3NSvrZqH4khhDH4tTV22tc1uO0N6H36s7y3tyJqiWl
XZ1M+rxi7tbXF8eQ7fjBq1X/YhmAOyEfguCyukaLIoKpQ8Lz1hRIFlxQ7Jf926M0YOSIF73mxXpF
uIcI7pHoaRwG5mHWRcuGzzESKdBI9qpD9QAadD1xxho5EuXWHGsh+pQh/oDtmnyg59r4lZ2Hlmjd
JQROate4LbbZkwWb7JGL/1WIQcPDyK5x1/iARrL/gJfAK0+0TmBexeC3eVG+yhQTNRsEOtCbZW1/
BwI5dePi+JAc4I/3vCl1HpgHnTkViHgvVNF1ckS0Nii0N9roynIk+vygz6r59yFmNQbkivf0U2IF
egkpWtZLjrbDhJ5lag10Dj3Vie9x0o4Clsmx57YR/Ma+vfJD3W5aLW+sb/DqLImD6CLsCsZNfwXx
MQ12OMcXK6DSity8x+ZsTM86HHaY12Vj2AyFJB0+1JO6INE6awiZqoNKxBFDqERbmVUxMZ9IpxzB
LusObWiDdWsJyHT9KRiCRPMjbJ48KiSM17VH9aDq7fNXqutA6TFICZMQWlOez3s7XyD5h2vLdW2L
jgMN6YBAxqdTU5Jcjq3soxkmascDOODf+eRYpMAGsF8kDMsC341fdVYgoC3McZolyjcetjEPofDh
yz4zigVf0Snd/yp9A4C9VYLuGhMs/ej+Z6b5is69Re+MrhAn1dR0rnEQENgbMe6dN1eFc/M59tlp
XxnEelL3SfZharSpcBgnvjv53Sk+LmL1Cmi5wcwTXM3xfHn5U6nZeFIDEDVCQR/LeuAv/N3ZiwOW
eTl7nzA3yN3GBaT3wy4sbUFCzvv34wfdC8x1e3zhSj18tdgv+CVfank9b77G1F9/Jlseu2ORbtxH
YVogJxjybZBlsd1P6nSNmxwr/lxm9WgqoDjPB9WQiDKbA165GnHKXzz5Vk9e63FFIewLtKTi31l5
S5TOY5GBg5plx+2NIm6WA+IWuiZrfn+wKUA8FK/k9aPb0r2eCJYCFs1u91hc0ghzuZ54APDBn0/x
LhgG4EHHxMlPbGcgzfxcKf/zJN4xNDmZEZVRdFsC/TuJ7ESw02Pn0TQdz/H467YQp0F0jTzwGAOD
oxfpI1LJp5uZaE3b0c9MjtVdZvQWU1qt4nYcs3RUZsZ12CybQZsn/YvL0BqY6ooZUdOt51oCu7qo
KZ0mv6oKLgys5ogHodgJCgdBwYMJTrUtGf3xJh+a1Ycr18I5SGJX6TDu1ZIXkN8PaRcZLQcwwlcP
vXn+ib71mzp1xrsp2AaC1Bg3OlYVsk273mfvxKr1NRsShy69KvmDyNlYn6h7pHsT054Enc/3SjTN
yMIYR8aRDL4IKF0BWhQkVPUgratH7Ipk2ak8vcRZqQmrvmqVBG3v/a30aIdxS53AYAjBxSlL1KEY
t2+cU35UZsO2CtyMpl/WbVar5bOutcDHxN/gAn3fuGxwzZHHpL1J2r2SPmsHhNExto+Pk9QI52E6
G++NdWGT0LlIqvWDoJvQz2ujYDN6wFdfZ1yZzA31KF7a/o67anfq0iHW2AFZzSR26Qv5Tir9aB1o
gTof2NHMxyF+ZtR1c2e7D0juaVgJ+jL/LVloWe2X+jmnZVrbtFUDifxYT4nymZnZOOPdVPWmxOkn
fjxk3be/RmBSWamkQYzG954rNDe/i2LITGmoa42b1CctAehhk+quvgy5/0ew6pqF6RXEk0mzAjja
qzYXSp3Ke4y6JAOpDstNOZApKei+UcbG1yleyNrbhlj+OULPavoLBVeyxZ7OsDPtfAFkxp3TytkR
4vjM5dJY2HI9ypQOv+d4ciLwT7wAiLr6QUsQP/GkxDoF+dmcCtu5TIRDJDezNZX0kSs9JEB0AIYj
wzIOeXcJJJ1618pVP/bIhlvey8JGojbpMIl7Nqj3vL6qr0bj/rF8FLs3TF/gka8q+ZDOEARUKGX+
BQOrEAcB5JOre7z2tt0BBo8ZbFkmbWvgiQk1k05xzkXhSuKd0lr/HnU3QOwfVk12RFyYbYyTB0JZ
pSNIlf3raRpV76/XhH7Fwv5tmfQi9SjX3OX10oRRLUCmHbWmfO+QBn+KmtAlECSZfQSkx0qSb5ag
T77Tn/F+FfD1Hp6+nc6+SteJ5wSapHJ1qokXwltgNNBAWVUVceQOlyYZHHSGRpFeLWMJ/E3lLaIj
tWvDjl/6iGAvZHqKQMKE61S4Bo5a4vtoegdSB3FPLSJ6LYsUmwNTN8mBtb8+fQRTTzRVRuNY/+wg
4g3VdBDWyws0i3eDdZF9AVCSuSGFUJdcUAtZz39G1jIdB0IKez9AjOMWCPTLAmCaTqau2FHxxOhQ
YhMLTwh4/k9z2rsOvjp3599VvQjQyzh8WB6rH1lK4Rw7LoDIxnWky0OdI4YyzEkYUfg2I88yGvpB
Qz+LOLZGHzHqYp+BySrx4kY5/mFX7FejRo5VZed/YpFcVR1eDMNm3N5DNXI/RJrZPAEUxvRGm/iK
cUwxllL7x09uzydoLBXhSj6tcGubBcXZrCG2tLlrFailkRNLun0TZDTAOFubXp+ojJsA3AkjW+yF
tTQKr5tLGTLdHNlG6qcH0z1Q/4U29Te9Glbk7vc1QY94ZainQEeHa4b8KDbYXoiDTMfuKlW5/Hns
UFRDEXeWCE5AvS/7mogHGDfXSS1YaugvoMdV/E9WHhNCxVePI2t62SVclAkbpXs7CnqUVCqlICqf
Xw7+Eq2rlv5nEjfm/U41v/+poM8WWWmLKOoZ2+Efn3DHiZxMQralxDgkbq0NOfmmMoTq+E074oOY
f368bNd0g3HNosRqlZ2Y/wF14PZIce1T/brmaOo4jTasxgjIm5xBGK1ZApo10i3iFeGkIoCXBRhz
7+yawUPMYawU6A3R3drZPpJqAdshLa2pI66eWNFp0a1nqV+2/3Fmezz5iADxMUChCyf0EyDxpmio
aQ8Aw8NNHfAMEI9rV+3jMh232Axo0BQ5dMLOul806h89JvQrjTafX3avZIaxQKZ29e1dHCkyYdds
9FwsTrsfIHtTzjAcRhqotQTSl7IDYow5XyvTtx5nzQFU71Mtu0CYiQfodABZ3kdxmVNUV6DR76bb
f7x/cWueLgyQTPKrCnvCeG2WnTClbVkz4vJtHdp4sx7lQsqgXjmo/38bQunD9AYohmH5zACFET9U
HEppKQSAosDL0nplpRDDMZlIn0gQD0aXdygcd9nIFRI57UgJnHcP7lHQVyLTMRUtTSI2vSd7ZV4v
TYcRBKu+kfiepwS9vCeQFBUanYck95U8PjMzCSSNEPplaN4ibm04tc9PIK1GchSbX8dupRZVXAtf
J6N0HGAvf32tOFr+BqvFQaUfWe8ClZ9eIInqD1kC7A7BY9b4LP10MRtsNMnX/c0DTGMxrJEAzd2b
1YlholKDjfVnzvz76c693o79FhMqIj0MWKBgr0yQ5MRSXQVh+6/p5CpcU3p2E343oiN0XuA4q5OW
GBCOsqXRxxZRsFwx+EWlPEWdsxpFlH+bSk4iHhcBbIISJbwBiyQWVz27E1dIBM7MyM0XoRR/fMhS
sTM1kxvYiz3R0ZEXGaUYtS8sWmxrIGan0PbLmNoL00n1co20Z+lAw0y3AiJUhGKF5WR27dUeKQWO
bwmWSRm1V9LZ5eLCGPe+j8MD53cEl+wN0DfdbP10s8RfFPaHsJkKB1sPKiVGkAtStyd3uNHxbZK6
x2qKVtOAhjkSb2Ns5dHB/M76sWjZEF/EFxQLaA0oAeWCz2SF3JZXH6rq5qylXJBsO3S+uYGYuNrR
nYhYICvIEjCcmq8lBwr3XyvI81GpGiw1ZziMTrixJ4YRXzaP7wgV9wfH4xH997uHm9pF5Vo7/hj6
dc/1OQdjybnViI5mfCADg5j9LYiZ9ubzcYYoloezVVGSkbVZ7/MK2b8YqZ6x0V81AwO6Ecf32AqZ
UF9iRqG6ELP4wzjNbfNSKKdLMe99f8YphGr6OOSKul8/R5Gn1+a5E/ZdfRmxsizAruKR9z+9JKgr
UdkaCm0mCUU7GVvIPF7bPKBQQzvmDf3TBqZf3H+scfJfXZU8RvrCJT2tT3hIeKBMYmpGfFNXyIBv
oqjGJIHeKceZ1ImdrFjsMwZh4zcI4Z3lGq9ItpXoAK5oNAE9RHcsOpT7Rlg8ZWfhukNBBm12wcQg
5YxG8YJ66YnwMeoMHItjdK/4S76SBpeLGa0lbtsgWFJ3b/vLRrk0CybQ+sSZ+5UpddWhDzYrGpo4
lg2xINmMQ0k5x/jjuinAH6yoATazVcs6pLXeUn+isi1/6vMxliEEl8QHEfzXZFa3H1d6RXdlmyMQ
tqeyGeJCty/Dbwt/erVY4Gu/ZBoCLEDg1F1poQUXUuG2gL51KAgP93WpisH4Uw60Cz/aII/dWsKX
JvwPyz2/g1d7LkgsUby48RiUBD1X0rHrp50uDLkbrtXumiWYvh5/7mB4f7BM9TJfTEsIxqzWhyXd
duqMThgc90vXEWMtkBIpE2ShdQLgLpqnULxlIX62fwB5YLt/+T5Br3EUy6B/NHJzRnyV583BtG7j
dxro3q2AWTk/ts1vrN3tObLMaA8EVi2D+c0IVB18DEN6hkn/0nftyMzHje0QksfWh1kHaU4FhKID
i9XdnSu1WRrn2ch/1GNDRt3AbHt7aPFkv+1wbn9eFVoQdCd3The65Mskc8q/KcSaCPUhOV9+l6b1
SKx+yKCByTkIsRTGgXebGdTP/XJTQgWFoCERVgrq8546scvumvNu1o8WbpDIfQozL9rzl3RrP+xY
GervUu+p0iYirSr6Rp+WN9k8XlV+Qn9MTpeu1CwmimmssrSeAQ+WE206wLE4z+ZikR3oK3JWvz4b
15Gy3oYFzmhzXG1J5QK+UXZ5ScheGxm5Nna9l8r/8quWLKjVoUM9+900joAi0KEfyRHaxj2T+NaZ
mHrD+j+sL59EAzwWKBmU8uMKiY37HPR7qRF1+DPfPNVz2e+mO3tWtq/gks/oLzluZGo95hfuuamz
KxlqMLeGeh8XRfPQJbv+s4I02cI+8VgtSTYWwjMXFiWJ0j5dA7RdDtUXGpBStw7EWulPsYVeaWOb
hT6a5WfyPSshUKenc4efz6vecqnkBCXNv/HLyjverjjALaFUSlE5RnIKbcnt1vPnTDMss+yNzWdu
tHn2fBn6KIhfKAp671fRRn48yRUGIlLYtF++qzLanowlNfZaGGkIYlxKt5+lsqsrTTwozdCVe97R
DWnyqIxKiMTnG/0aDAOZbleD66vtVTDCSB6QtFmo2O5DSZzgCIALHvF+m14KvaqPtncQhoGn2usb
tcBGj0kTrKDFNYUW2nMSfIwgpj+yg5q1YWobg5XJvzRkryrRMc/iT44CfIvzy150tv+zrK29XC43
zdqduYwyRtVAmdipnyU2RCKZCcY4OfGEDHk03Jkez1P9rFA1Z8bS41BsSy0F1tTLv1xFr7u8ZM74
wSjx8T3Lf5ehNQ+aXtOywRLbhN1UN5dWrSB+S0yWGFsUJ9c+cSvt/l7Yjoy4xv0X1Vy5gAhGl7dU
o/5h9JkVRCOxMjeAeqk/zCqlTHl8afkLI6Z2jlp/Gnb+l8qMMQCuGaMPxISpBEXNQWBSfRyriMwB
/ebD9Iq3evuCqghZqJcAAbcfHl0wOaD9+jkZGj93QTETtCNjPEjLtYxEzskPq0/Y9Y/jp7yJUIBg
HgHxghBfr+cjStn6RWONc3lNaDkckqcBckzMGdqTBdbNkEk4qX/6gCcVsIKhxOllHUmfbjoHt2TI
zUEcsK6ygE29GPpdp3z7tkhsqtiDxdrhxlFVaED9zaM52c6VO17POmOhktUCelROgxadI3V3R0EU
JjL6lAjCPMJPFoRP5QnRIntPzpIlhO3uYe0YCSnh27p+VOhnJRAF7bSgi26guU/OvoVKYOCjIRaX
VNFw4svZz5eu+++nyDn6WciPVNBfiRN5UfIX8bR9ilmWtRXp0wncHUX+fBDvnlOiNVb4hd0ar/Ce
9WXFngCLjTETgDGiVfvsH/+3QsQS6SLjKOQp3H4cM3K92Wq8aprag2uE7/VNA0B4WMg7GOgy7Z1J
C7vPCJ5nrMNHXyDamZKAvUVfZx+mx9suFOYJiSVKZDsqFWkRgN63PPYL4rjWwPsEaiN4xPu4NQq0
sRbqrGZV15pyNbqDlmbswzEGxko9TR62+gmEZx0F6yEzVZtYLSUrf9AowUGNNJlpRlvv8sLwAZ+X
N/PyqsA04jL7By+FykI89zLEtdi40rkqcZmsssblO05WOSsbgfqxK9u7Sku0MOWFKoyiBeH5fHo+
5U26P7+JtlYaysoC/xzWVB+xpxOQaTf9f4iQVfiMadPLiupqJpM8MCVO4zIAJXa6NL/nBMKQYOO+
RxXYFrszN0fHySe7XA/rbcIkxuMemezkT4Ms6waDLYAEUkj4p2jpiy1BE2HkPlT6jBxwpiUomHTv
0+YniB3LkpKPsPqFiV+7yBQHi9hBM7DbapA1ADKbF+MI55mSRqB2QbEMm9OF5FQ3f/PvINsRXfhq
vUSRStSZ6DlY41xNWd7vH236FiY9Bg8ku+pL25yv4pMOuuKHFPbpWFlXpbZ++ZLBuCWtHzxdHQgZ
AWchmnm9RHnQ9wTI5XL1FyR7DDZupliCbDgx3Q9PG6GLDZq6VQy/XzCEYQonN9LoZumCiz5TLzoq
9YwdPkxdHf+qb2CDXJ4F2F8n9UvyIVEoF+ztyhecLGkMy/IAqYitAjK7lGAQGMeU8Mglw1x0ifnX
zbio4YsdoYVNQlfDB9onGP5JFpH3xhMoHYPc7FFnjzL1haHyvm7KlJ14s4RZMUbJZ9DTumNwqMBu
tamCX1p0cGzJCNdzIyh6pSFWvksUT8qlnYh85IbfKKvOGGUQzPlpyEPH1LugIDofet361AADTvrx
nLhkic+iQYWDXcE2OQRZmDHp8oWm5wo6QtovPlAgLXS5NVoqrb0CjAUMSe16YFmglI41B4Fc7ybx
8PVZqzppG5FO3XpwsdduW0ZCMOpx7pVH91+4YhZ+ZhoLNPpys66jsF6X+V6xD8CJOFc8H1frLsu6
gfpnWfUCcsm3s5tZAzDDd6tpk3kzl1efu4lldtuBjsi78F2pTsHV86MkUnoyM2lmA3nYKs6nLkTb
gCuo1WJ4OsfDNXSodrQoTkm1WHKxRXJx4CyR+OG9g3FujqtFfUlGHcmj0mjQhwEAb7kf54waHl5/
yviOyixJxgtKf9ibnkRHiHwWt51/v7DN4QRZXTIkotxRByawPaQgwFEdcc2+VR9AjG9anLzdGslg
QICSbZX+hMjWgtLeeb1QFk7d+FC5EDouDWvNrDZe2AzxQDwkscyhyVds7kmKEu+pQKaKwTtWVKnI
liTW8qGMhcK0bGgTxGRtXGp2g1cJanoQKfgsNRR0xwoeX09IAAg4uX9bVg4M3HC9FfAjFtxx6CWv
CR0pC+nKxoLuAbhpsxdD2W/4pHE5IlNSwpJLTS7b8o62ssIwdB202BDDmZbQeg4+T2gfTqtCtih9
wnQy/NhxAM5D39zN6tzw9Ev0MPgJj18wyguOeJhF2nCkXE6ARYt0EzQQ0YPEvbN5fs2WXmjNR2w5
Hyvw9ytmf4Xkx7v5f1umwAupJELwciZtje37ENctbD9eyUVjwum65r25Ql21wMmfX/gKEZaknPS2
jQFOKuChRVZ1CC7TBThxrhhWS3hY2LEW3Gcrwpg2jaKeOWDJSDVlQ2Cd7KmfLya0lDlOO6YTV5bu
FHEdDRgNfRxHb2Q7bqNVbykCu3qbW/Ri9o9buz98uykCm83OOLFkVB8i87sedrmg9n1B9sJRdUXO
mj+Sa6UUOJ+gPF/J9cXgLOiJM49PAM76X6VOSPKCAI2czofkBK4lWhSDggLWvO1A88XCnp9IwTit
/b4kNTTVB9b+MvmwFgRhtztdoI/StuOSrLfqGjbl+yGhiv7tr5hoC5p3mxI78JqFFrX9P96GcLv6
XP3LcmxIir60zSFaXVyIifmrltvRrWtkisjDFzy+FBvK4vnFZVZPjrv+dKC4KK3xMGyDJS5gW76W
IsPUedca4D00NNdCIkcb6WvRqGpElKBeOjiZJv4xsZUsGBtirZdssc5kC3wZhWaeUrjw5+1NQpcK
98zv0sEq0RrRkeiQas2lFRmBJ4SPPilH9IAGnHcs7z327ZkkZQvFNd8b5TNXsQxswp5ND/Fgo/bz
HgxbujgU1xurGMZvL6xlVFs6AsF9TdpraNi7kjlONfoVYCd6sAtxcuszLNnGg43ImhLSupwa8mwe
PN4ATLl0C9zV2cyb7e2yZySJtfWGxNRfqJ8HloFo7BXfLMghbOgZOCO7X2ma+vAynR14bsCgPxji
mE3Uwy1J0zCtmp9r2NBE86rFkts9/iouoWmTIuD7JBZDClLBLd2SIoTFCDvMzI00kt9RC6wDObmk
uDRLOzGGW8wLBVAdm72uQH9AAjGBJzSWE75dCq5Rz0jtRTIu3zlkQtVkm17vz1Q5v7iOAIkWBdV4
QsFHhfzsBPgpN/A43irr4mRO6oNMIErjDB8QNQwjC5Mst/GEXGvaU6X46CjbR8SjGp25lKTrRa3j
FtVZcI2uQLk2XHNRT42zHf9BNWPOmzJCqo3/FTRk1aR1YRzqqz6hwNPiCW/mO7K+QPYAeYT6Ncn8
7aR00or4w2I42DzxnITNQP8NtzN7CBY8uNoIEkWaGwIiDL4OdlxMmL/GaKTTaXKL9m0XE+vYzYK/
wLnEnXyQXKIyMSkzB4c04ReajARPbGVyYsgBgyj5lt4vWdq7JaxGISIyepi/rKgVnwMbS7maUEj1
VwThbKUGWQagIeKDgjfeVHOdKSFQ8kn95i0nQvpuxDgEjseIhAOiQPF5/MHyezogdNMVjMDTDi6s
MRjW1G5xJX3nGjVJ80LNg6XkzgCSvHe6hgr3nIcWo2NFbbd75GHYjFoKr18NFL8tvkYKQXPa9cqY
oFQROOWNVVxOTXQsG9k4LDSQe9PYroNK7SrC3PVptv1wiPcEPGpfCXMHO/arSTvQLyOXVQVjUg8Q
94CSMkH0cuenIuR2xASot098jhS6XRMwhFfJDtyA+guB1kmko4bUwRapUq4bw/uSNF8qb4k7avPz
5sY7WW3Vt4fvbPAUdke0wfZhmHfQsKBaR7ZSWBZjs2qmffVWj4aiaGSMCEjBCegSKJTjHqJhgtFm
piEKBNd1scrZY11b/vTLD9CLoypbtPwpNd+T62YYOE4LlW5RjHEi/PpucLC4O+DAt7Q2GeFgRQ7M
SpgFo2I0H9aWUoasOHh9WJFr7ebSy5n6A0+TSWCceej7s3aRAKCyF7kBC5VE63oNnWelseBLUzow
HFQvwZ5T5DGH11hlpgxSjNMtBZr6wpF9El122/5GDes2kQyPDpJYWmEflO92loGE7XNDn9R9zoGH
wBpMabqsPakWWqp53RCdroIziHAs76zg05Ci60UmjEuucJ4kHMbzHmmU5HyFqJRDIAG5C6dFZb5Z
uF7O9GGsojbiO2PQNXbtBZhKTRsV/aUIa45TZJcWs6JERQBes6xKTCEtRAKV1za5MLsJPt2PNJHX
cqChHmIE/xYqHf95b1pBpw7Xd/6CLmGx+ubTUMcoptqDq7EB6rDith4vbThYT2k6IooAngpeJobu
MhairmHT04Gd68hkK7mwCrwrE3KeBVLE1y+jz81yji/BiYL0lG8ehj0Tyy+7jpNsvUNL1AEKYxLH
HieI8OF1qCbe1MzGWkZitj9Hz3IQJHQEx4brWGRWqZHGLJUY7T0gVPzT1Tvo7WTc3ziaXns8Rd22
ZQJEJ/NiUdZZIacvJouQQKPUc9ODuD8oeDt/Gpq8HdmjOUANTsQPSHSStsjkN6isdFhyfF7QbN2O
xAY7hMcVewd5CZNhET3xQOuMMc/1LAfA/Os2mSreTtkGhlFXYTd3cnTDGI/Ppm+8ReCekpX44TvI
RVS7OU4AQ8SfiMuxCBHgZosE96Ochav9Krm2T7TAQHUUbDVEGIaeYmKihiqC7wcVrPNEthEXWAV1
uylQtA6/vSUx0isMQcBT6Xv2olztn65DysfGrWaul/dWbcaLha0eaEgW/qDTp14/6IZ3QaeFRaiA
hAyTvHvAw0NtirSeXJR5dotTitC7kYN1djSNlVu5RPrMTFbEM/zcFz6Wm0ZGAIa8gj2cki2dAIAK
g16ArD5BXwwA2dDjiMmoz/ylLySEdCKO0pm7t4FAUyQQAQ/gjfi5GhnWpqmI4SodYyOSUY6Uuo7U
aEtLTAA++47nEbqNEfgJCjkhM3sZntiUSSZ/5FtBvrRqK8v/oeT18G1b4CI+qvG4obxkLKVcKDZF
JnxgKWXQLJ0UBrTU32BpeAnLpUMaeDUKai6ZAIL8m9x/DLEa9CwA8Vmr322dLS0oY9gxWWZvjNN1
nWQbHJtcWErYdHX5qKFsV5XvHalwV7Q1WWRORvwAoykGNBMryEWZoYNGaEcVwwRD/Qo+acrVi/kE
qPfnEtVQZAgIni4275XMfhUfMwPsnPYmxm0yPjeanZHLB5YzA/YJLguxdMj+sRU5y4eD9SgTHo8Y
M3Km4xWgl+vEfgQRLVWD6QT+g9LIKYdkcBVPB5rQb03v1x0CTLuusr3f7hlidUJ7mVHtNKpiXJnZ
obkzdPstcesu8bkUKJmORMLY9Ki1nWs2NK3s5151I3L0czPUjDi8FPJ/fxmEt6WLAZiHLwRYyRmD
v5yX2ddPkVXhsXT386YGjnZiQ6R62ztCJ6+YfI+x2HF2aknHo/+RUmcmE9nO2EbeJxCDcpevLLwb
rai6OQPV9gYa5yCDqG4+fcrMV+RgZ2HnsBstswWkB+32Ge16r2rc2mtu2O4pRUnsr07ul0gS1A3U
lSf6gtfeu9YuhU8RSY7g+0rne0Gmt2O+d9Tcwcq1FVtoEIEjuWjK+xyK2saEqRDN2ur3WTiQJv1h
jPyAKd7VOoeM7smWnzHNs1wlS7PlagBTZ7CrY5cUflUAnYI9QBcafcDs4IO6aw3TNhceBpynNduC
MvNgevgV/pQdQis/ZN9QsKwtBldoFoCODhr9oWob1xhxgvJnSflSbgpn82R9AaWxWq5UtR3scDTJ
Z63iB6DNPrkLb3T/SV3mhF5k3KmI6pqknPgnl/h7/fnHnlh/oINk2jyI9BpGnunkg48fvVUMXUkd
zGc1LjKDHqgXn5iqO2fjMs27sZBWwxRjeSl4C+Cabqt+cmmHMM7Tswq7N7I03sludUaf87lCAABB
W7tyinwPFgRh2SEJf/rQ7eqwg6IKvLxsqA5YzEAf8MAHFKPqEhWejChpSATUzbgoL7v1aMXmy2Ck
pC0t0JGZeeRsUF5Yk50lm8ufbZLjUh/kPzxwRiOGqPpePB69a4k67QhqlMIr4aVDTUZmE2Idz2J0
0Lu3CO0uKHp7ObY1wV1zKuCxN5zCfwWWod19gbghMvdOQwvDKf26s09v7UF0W2Rj3EE9B8I0i6/h
Qt7yCdO1J96XvgZhamn7R1yUYhUvA8SEDdYw7BU5dT149/12TVSJftqD8Smcuq6+gN+ENzzpjTSr
1DUlTfmQ8v+qu7sNKp+zbgrvxkLdJ0hqUr6NusuDvUdzrcPoHIOu+vzojY9cQNdQBAjEezDJ33Zk
/NLbidKlQdtFJajSyx7u+JcgTtoCDodPRP9uRub4ktHp/OVYAk5MqeB7BQph4OENwpamaq5nYT7i
3FVShoEvDGlp62n9pjbgSA0eXh3GyAP0y70Z7wPlKLwY10irIrKNTTVHxvc/hz7amfvO3XXK9UAY
IARKVNCZSHPXPQAz0EEj/KY/0YwHvCHAUs53ftz+9EgGDstSTQn09ahLpdOYS9BX3+OjFet9xPnK
Xgvo/GYX98L6oHTxvbTSNmvnf0WKgc1MqGF8rFQIHLLLL8wSgzTHI4eYB8oXBaIZQ1V4Yahvcusw
FhIHRbze8ool75YfLJX1pwtCOyak+dwz9tb+a6WNaqJdmoZefKBNojd91RdhBwQjfy1VNIs//Xu4
L2u+n4fUmnBgt95HuL7N1ATvpRF/HisAho7BYrVTuqR2JYWZpcQLfkQ7TcmK3BNoa43BlxsfKF78
gavetWdzjsMd8iUiu60KPyB/+qjYdPUapv9w3FhlhQQQQd3JRuBrl6Upm04qkLS0ey9NIw1TU6Kl
wTpFj4ibQuk8CrhTU/rLByR/pLe4c/oZ+EU/V/zZtrj3c1nXdrFWJ5V3I/NkmUPa2MSzzt1q6Gf9
7FfOpbLk4c9E2QsshVnxbO/2yEs+h3q5M+cQOZ0C9b+f2q87xnMrFqm2PC0qpA0byQfAOio2We+T
Fvpk741iv87FeNkVlprmBXIficSagTV6wegv++Uw39KT09zs0aDwkh+tfHBjmR+jE33sDCwnhGUt
G48Uuc6dGE6qcnnT5fyFlVWg9q1214xTQpqhwEaKL85BLOHcrwjC+O0oXQddraRDNm9pICkx+kjL
EVWis2salN9tLcoOuPLqv5mV4H81Hlw5IJK0dWwCe3sLECyT722YfRlZiFMeEE1sfDXVpsZw5oWw
rCgZiYStSEylL+6SAG++orNn73yFKaSLMoDVUjHochNJhs/NNNzqtyMFJcl38/+68tIO655SRyPA
sh3RzmpCxlLbwv575wFfkFecC891ohkj8lWDOxH4m2e0RtiaJidBuuoBGZABh+/aTkRAcvUkAagT
8gzeWPWUVzjYFOamiav/mK4iCGTZfFQc3LCWadKyAypkQFPOv1ShQyHUURA8WZknIUyWNjlTPhMT
OCArVP5B/BIFaDzZQ3iWGo7rp8QhtVFxuOyPq4uc6VV5aohg/xOAJ4fcDy8/GPLIjU5lAwgTFRlu
wVLdHbCmWDJciKyhHimQsWWMIxR0HwYjSD71LTtauhL9a0edYiIZ8OClv1woSZ8IFmHXwxbn71TW
2Q+mDJls3ljEYg/lQ9h8ke+M3sWplaVp4lCEKxxdZsHlbG/lIm65OIPSLnYmfncgoWH8b9rtbPll
yDkYyFUb4q7mgsSiq0xYfPf3524jrreJME2TpMcEIklgZZljYArvqzNamnGnICcPm1r8U5msmXaj
DksrcHFY5mrw9MXx8mppElGAGIWMR/e5vwMyKA8RXAwh5cgTZaKdI/93AcsYYETwjNQAxqiIcaYq
NwSs07yO6f8eLfn/tBg9faUljXNN6T34z1zBvV+okFXfjzdiYrkIBdVfmsQ7j9HnRFbHPkaahmEe
kcrjgHpuWJjPG92+GQ/vi/RXeRLNg8RnRtGgZ5iBXc1RImN3YrJn5kWUapnBvuMlQY02+Sj/fSeN
AUdTjLLPzTI6ERnQHJ6J7lYkbqfAeZ037+/E171XLKYeGw0TL7F2MYrWdA/qVxC0+wVEUWZIEV01
mWJAssGgiS3NS+xp6/3wtdoydRKJlEcsfdaBYJVOEq1GIKwxQREAAcNiHE9khtcJEj8FCRehh+S+
YFBDlxK56PmZeDrDidg03rbGPdSKXmtGQyDTFRO6EWL6a/YdrIkWQjGW+akpPc5niWAax2KMymhW
YOoAj2XWjH/ok9iIAUHB1Qvi9EMjdSMJNyWtKksLpDS2PJST+T+l7UCEe4xMYEQSBfMJg1BbKz9u
EfxsT5bn6hGY3ddcleAZ+8u+Sdr7h+hRQtyCe/lgdxiwoQ8H0PHVZp9GY+0tUGhDCow3s96I3fXU
oXX4R0jTi7+896UKhUPQnPuTkxfidlBOTaXwB+fk+QLjMbmsW1P2jqVrUjZicbW6nYL+QhoJoUOP
uwBJQxI4bYzWJgU3hrzNWZWPHKgD0ND6Rlf5rHTRohhjbYPZ//FxjvkSfSA+pvYPJTllEAPuTZbH
/sIjaPNapRWAsezr0ierTmcD/gWAQPD0YkUA0jNijncDURw7fPI5UzthrZ8DrNriPEHl8Jx7mdoB
8J+I9yvhWFwkmixX/McCJjE/CKFHaHzDvhdWW0XhIXuxhA3qhIWilG6xJE6tcJpVcz64iJbP8S2a
tCxr26Cz4lNSg0IRciyzV9/P8ke424413Z0Amt5aHRkmCRY+5NsFr8D6kJfPsIgUYTUEPPi/L8cC
RdN2oMj1R3QPBsHwq4LiKWEHslx3ljTUZz7YIvae3xpwNL6E/9HUgPRaV4x/VjzJTfIsTPQn14Zk
iqEd28GnW8OPA9n+XrbD1DRIlxwgyR0GcZrAT6JLZREXjr4efexrmepdBm9Lqqka3zp1BpdzySKm
p5kEflwWyjh773lz3+mY4+e9aAWRsb2LLAYJiwo+8CDEmUiWEVhr4VCTV3s3kDJU5+WJehldLlQw
YCD7ne7kql64jzYfZIIcn/O5Yvr4TAIYYY5Wtl6jlynDH1KWHAxA/DqeCcqEPG0tzfnsGe8PzWI4
qkx5tSm5+e0vNuoMit/PIcHtI/RqPj7UnzswTXUEt/TwMxE7iDQJCZO11Eky32CZEMJL48tiiBjZ
dgQM5eRw0j8eKi2pVvkjPhauz97FRcQ+xuYQJfYZ3hICxZLZ5zbw99sCvATj7bFH+pB/REOKCwZj
FU/oOx9+EaprNQdW9Kwia8bDl02UupymHZ828i03DV+917lbbFvynJMQ7ua2qtz2r99yuJ1mecT2
/zTuUBBmY0sBW+0Sd+7Efp5xgvD64mEw2RadxXzi4M6fnrcN77xXlBWpEMu7cGhS5phNFeUL95lS
qwSzaqIvQz4xlPWI0Yl46imMEYHIfGWsFoK0aTlQfjAmZXZ3m7TOjAp4tJgO+aE5MkGRPgy8jGS4
17JqrLrdVHpdcYgaA2Te51qJkzO6v0EmZ/wWqMfQyn/naNkUxiOQj4RjtDIx1jH2tUuXqJqDjbjs
jjIhNwiABVjWc04/Put+AOZLzan9WspVw3SmMb8sOj+dLgPlHcEoTlge98jmwUZMM9gBhtfOmSLE
iqHbiPYEhFw/EsV14auWAhzrDKvv6Ck+21aBNdVZl12lP+KQQmVSN5ZQnc5UXcxBY8jDp18zzjZd
8TnG/qbo4f8ybO49vg0PP9oBjcH+0ALMpcjfP8j7kGKMeOKJRnV1o76hZPYDVf1/AWEAGzyAlLu0
noo19KnibcEKS2gaUO3XfrqEwUQNPBBm1F8+1t1mQEO7CWgpJWuaM1sSb6zjabgKBm4qZ+s459CY
6Gj5iMSctbfSquA9m6qLaASPDWSyd+pXVZGT2CsAvi65io0I5dJlP/J+WDvHO+ILI3VT13pDXzOC
8nx85o9WvdlzoU1pcpiqUbWj0rWw8wrHL05JWLrGxdLL0DARloisz5K9ksMAjGrGDySJSAsXs40u
ex8FEp/bj2G/DMcFBkgNAupP8ABNrIdV/l8/xu6g460JPktyM5CD119jrGC82pPmRJ9CLBKojpTU
tngM2CBZPUpC4Qtzn0Na8JjtVct5auvz7Wf2cuxpv0+ip/fV4D431GA9dqIIcXmoSmdG/iRwtR89
awuvgPEGGZXx4gzvpIBwX2SFaPjF1mIE7ivzQtxq2OyYPYQbdvw8Az+Tx6XEvP5XqTgjKVqhzrOQ
PsA/e7oshBeYuMBssoN9XBIjLKxDBhoqkPomjiaHXqw6rZryyAZLTp20lOf+L7nqqkbIFR0Z4kVj
R7bzvQra9rgaugqFWOEFvsMrKCHtm4fBGPXs6yfOQR5bL0ELJGf6MbohJmldgEk1HbXDE7IiIcx9
EZAF578ZJuPHkv/gOHl27kxJPLq48xGKz2Tri9mxfEOvr+VdFL8hX+LWRon6wS6Ku4IBUeEr+s1S
N5n//OYD9VABct8c+fTnVmrZBrXs96UwddX+u/dJtUm3G06EK3at0IzX+VJn9GdkE8qeJAWcLwWo
2ZhgiMOqWB0kjbh2/4dt1I3qkTCLNw8EoDAe+O7UTmquO0NP49hU8C1U2XF0MldrGY84rdY63N1H
E9F/LSvmG4xSHNNEn6iF6Uaxx/PSDm3t0q2hQNnEjP6z3TsxXN/g2DkKf01iCZpkugDlkSMrqS2T
iJn3pd7YAYDKvMTCU745K7cdRnMQMrCmiD7gKOTjLVME6lOzRVTOQQvFe3M1IYmbfcvXa8QbVIQg
s4X+ZCHnxHEzDHF6bCbJ1wqVjLJT4U7zP4AdmWjf/LC58Ei8PK/938TTwuTvaDCq3VMpahJG9b3Y
s5iSFICB5X33QLcpwu9G5Q0wYYP7LQJjWPKygnZoFK4hgevh8XnE27ju/jDJa4V7d0HF/E8x0kLW
Ei0VLoMvjepFGHCsqvCP5N4d0trvhI1AKLiZJz/YN3lJ0jh4fEMsS+D0cwBAyH2X2DTo5HkD+doR
rj9TEMFMysL8u21KZKN27CGaFISfvadEUwfZg8an3BYb1Fw29XlOQdZNlrqgp6tyvtXJE1v//E2C
FAj0ZFl5sytJEgHIth00soDN6unL6RJzmk2tm1B5UDpQE3GWR+NhWsPWCrS5CbYJB0SbYwjRtYYG
1+xXsVMvbFX89GacN0s1wZqfy2uF7N32uv8LoFZpd24b0AcoDT+uWlN0aGSkL5oOTpXhT0AEkwhs
qDCaYFTPocFnLEj0fQf7usRO9T3egO/3qdzTUQIMo2pLKmRNmUmY5vU51iWKwNnlNXyX6C7wlDMF
Y7AQbipo9eM/9Z5MVAW1JqSszg/bk0zbTBpzApWYaXCNSXhFOgSN2hnYy7M/hkcnbHkNyNxag8nn
hTwKm+LDZMOwnEhrUx4eSDZH0GEKXGaSglPgIjj3stSH2NkI1odLcyCS27Ru2ryjnZKhuw+PayCp
hwiDRQUQG/0weieFkb00fZ968P5/0KZKyd325hVIgJ4okdPYno4svFFHOuEXCFwlz66ahnIcn6Jg
aHxD3mGy6Tj6iWqGAbhXc++NDDoQ0x3eODAMbimj63wXLOHU1qxTBOXr7iqRzbN17qw+5mV2p3mE
LBgRi20Cg1bCAjfuZZVxTFtB+rYGuiD5oU8CdM1mCX/6B285+6s3/WKkpmzazBERn+dBVMkhh6Ub
UfHuUCH5v+jaVdUUVvP++Mk0TRb3bzGxj3xYXA5nxYryYtuUy56bqi8lYiD4RG5YE5/PRp7K9MEo
L/A41SZcHMWN8nIH02p5C894jp08xiBEYxVGjXyswss6XRE6V7rX5M3rKUXsprByu7kfogD9FAOw
FlAKyEF2g57ihF/9/xRfAVwrEggNNs+Fs0si2Lx4Fef6wXdFC75X0bAFCyOb3yw1z+0NzbslKL7W
OPMC0vGne4CJ9eh/pS5oiP6t2OHNuViKCALXtYs5a3aWvmMYja4Ds4XDpn2En4kxrNdNKPceEKEE
LtQ6RlqLjTIA7nzKQnp05SgRQzeNd28rqGdgnUqJhJ6zLXrTbMCe7wDnUEH6UwoLAX91fgoVugcp
fERftPkef5PqAMJxOxuMpizH+zKs1CZanQkEErX11hsmAHTF3+wKcTT1y+eR898hjjm+Tk4+vDry
7xfNi0DYRQuh4zrDgDjbRKRMuPSDwEKzxYBTRQXTlY1yqJqzf3HVCkc8gnSjMNYDEuJ65EdUehrk
C7q7GtrFgw4gB8zOzQpERgNQVcX35xgxTiLhqnG1+FhfADHZ8i1b+rlt+PE+lQkaIgS3IAoI6VOY
ZEmyzJgphPwfmevlI2ZKOdZkhdYPXFRQvwcmNMAye8avXkncdc/oz2ulryr1D77pPv034yz/XVY0
CbZPBIKFj+yVZgi9dFUjgSuRrTDo9n7GtZFBTeYBmoXxrCos9oNzBfB9gYQ2y55gmwW6/kIiIK1p
vFlEfZASy78eKtQzAJwk4Bv33dq8DuXaDnynhEya0tuYyk3DpRVPtULL7YIJAFNgvSG3T1cxSjbN
C1GbZgKyhxkqXsyC/9qyRG5sw+ba/6AK6tqTAGsgX2lBiE2Vu5mwzbVPZqGjqt43dP6I0XcOYRbQ
j1GRT3Eh+/wzBb+TTge5mVxS3B/bbMMZkg7D02HRCSwUXTDwfGaEcVC/59G0uIRHLkkt36kPot/D
1KFCrQ+0GQKXEZaJA8vL0+DwTHFhaiNHt6Tw0BlpidFNBQpKZvugGuS6lqN/q3w12LxDsgs8TN3E
zoaIvDqQom9lsDt+TTCf9rBxg1enmGWntAzxIVeVOvpR7OCAGRmvjXJ2okmE47oFfdSgfYbRiNKo
VCFPz/JOF2EX5eN9SVrarx7/UBZKsvg2pS0Y8YtlIoFXWO9Of5TMDojxRZqZUSErM+Q7HYKqKPq4
9z6v4/XlPu7zjx8CbIcje6Vr2w/2oBuMzizlZzc238Ari3/UpRps8AYxsOoIVirglHoyrHbSxtl+
SEDmUA+AQrzdd3sEhI9uHtraqSFu1Y6A2YS5RmSmpyNb0l/afzBQZSXAE7dXi1ULDr6CzBsmp+m6
xwO5MRZnYLn/zIlQIp+JeHtZvhCTVQNgq6kjp8wbmNxGCSD9+E3UnKp+u7tfMy1U3lX3hfGDJmDu
UPqNXp+/YSGeXInDf5pYQ1n34irpr3781PWz8fz3MvkxgtzpSD1RyObQ7ERo5ELFyeJZx0XGymF7
ZoAnK47nLjAPl4B4vnXtAZ9Q2brHTH/RQ8NY97vbzvIDNxRUOeFAqGl8B89mPPNGxRZ/RBEl9LHs
tvj4UxkScBgvzrAT03n4L6yChB4lFDKnM37I4Ycijw5lM8YqxzuctrdAgBBtRKdsfaVSDHcp+xq7
zG2fN+CRr5HqOH0rf4v04na82mVgqn1fXN1EzU4sGMSCilrsWczguscMuBUI8S+5wdZvJv2tMgN2
MUFSlOER4+KtR8Z5Rp5lhMv3IXowPCpqNYU4Sx4imVBuJEHTfGEjgSKzj2chObltrGbOeh46yMzJ
maSm/vC5xQDySLsEWTpkYRtzIabO6UFEMLPV/RhnQFJuGslQU88xRxVR4gCVFa36CUY/4btxmASG
Kt1UGZtyXf/5PI23xQ/il2TsW1lhgW8H497fCCMITy37+8rB2ZKN4OLjuTzAeobLqHQcMTx+YuD1
0OYn/1CXRVba3vhswvk44jJyTLarGd0fNYSc+N7iMIlLIAc+CdOAuMEeIcVv7Romv+5kTYGDMWM6
x8RIBav5luZnWokHCZ1Lxkzqd+cPvvyB2ZsV5xSc/PZ3aREBBC9bFA5EVSqtBCRm+CFe4mFieweC
AyYOxcQu4O+Qkd+oPH+pQKtax5aIh1vcdJOPVoAwV9WOJClx5ZKLxHpIhGcgURnrIpmGtHQQx40S
HEXlbtKP4X3JeHrolIfJQ+KZQsEHc/8lSyRpB+POtEp04yl+vXb2bfZLHQLo/MxlQWo8ycYkuwj7
SeeAkvbNEkiFwbAcnRBpKtTKpD2ZaQ/mXroMt2Bdm86KXPM5D3krp/qSlfBJLkKLzIHt/fTSBJuB
9cowsLZLIH3pEkOy3rd0Jgs+tLsQyMltQeDEmb7x1p4vC+N6lCRioRIZuymQYUvm+ZoiKdksLYe6
qUymXAjYdAwtYYxEawLYYPdMfASqixgDT7hXeMoc7fAi2BGAv1lXEqlgFIaXMNkUsCIpflkCilOb
el9gx/QD7E+60eAcmIXT4GmJtLvBeBjU6KR2ga3h5bXlHv5zOpKlZQYgCO+EN8WkW1nXzDHhM1do
5FdjUHXWM9M7juiA2egjekDKsMuPAII5mzB4FHEe8vnHLUftEFh4WCTRHSVw1dhMITOHG7mNvW51
qf1Nw59jTRuwgbA7WVpvg5kcGSHaoMWlSSnhIFwiO1lwGMgLlOIXx5CXZo1vAAtyFyXTvruNggXf
vg0/iRjiGjLGHMCU/YLpYsWdfBrd3wETWuFo7507ZVSYsZwqq0NZLYOf0Rwe1r5FCZG3q/r31zjb
HkMa52AyiocodkpYX7u4853IE9XYBWZThZLFUdVjKAgofrRgvQuVZA5ivUq2R+lMQcSq5EcSMXyz
hrAexts/lw4mGuPy8SjwrI129ME1U521xY5+na2Oc17DCx/meSAqN0wgdfaeOS0mlkrg4wBC/K8/
cgKnq6SX/Qk1kLAYNLPXTOhnQiFUZRQdXkZgBJ9KRevvw8VSSswXmpFNx2FqPyLnndQMZTrI5Kb+
kQk66n3psebF81f/yD+tZ3qrkza6jS84R9oILgww4kwj7q4iyOvM3uTtc2jVKWUgfvOtFE0+sSY4
Ro9w423gHS+i/x+A0EX00CKLnghAP54n2BO3KF9mefxNUsg7tnDDJZX9IqeZjOwWyroKcyHvxGTe
Lf9yQuzoDMTpYmQkxQNrVaMDI0tS4EjeHEuezczV0RT0dDQWcSU+G7eE1KEQZBo3s9b78KtDL9CQ
vnJSHYHrQUjAgwZyEJuSySceMOvH4dWqSyXun8o073UaXag2LD+lTiQe3OSxM4RhhkgVBdJ/KkKy
tCdlpynjj/R73fa51W6fEWsKzDpuX7YUIvOjzzqm0cuPaDoXvTo7ccfmI8VwTTSSSG0PxnBeA5Ry
hr85Q7O9svlTJANnsJSQQnj2BSruxOHkStpthwvmFqUUh74UMi5CGgG4xubPZh9q0BJOX8oMSgqI
DsBKjoWiKyaRAo4Efvt6cVYIBJbTuJbDtKBvUu7/fmW6IqBDCxK2LFRVvZP1rf+n/YfKaSMMfTjf
n7Ax5u76KB8Zbs5HBbmnh3bue37h+umHCXckgrOvpuQShaVKcjbkrsK9EkVpU4Bsbf4LYks3zrfV
HA6Q6KkM0NItMEWGyBTrTD56ZBAjkxB5biqAR0l88RQc9WhGiCJuf07fRATt/nrxDPvKxLOkWu+k
mbYQ+OA99POWZSWKrbIyWk4ohMTiDHKA4USzI2pHEaYWwj/ixmPkJRw34IMScBq1EbcA0pQlu63U
pmuVXiRw1nWI2GdAbBhW/AiETNKznJxykJ7WHeUKo4MTpljLzfnihvFp28S5k/t2RIoSzotFs+si
4rsHIe8tocB6Ge/FVgP3jkuub5ykpZineBFq8b36iMRkJYXJNnGHPupaLz7bhYJ80a0Qk7bc0tVr
3lg9Dd1CLwwc20Gm0Of5VQMjjGPyhGshJ3y7w8BCwx23+uT/iKLyjpXrt6LQEzW5uDw0Q86kjJwQ
vSgNUsr3gFsp2u1k5pVlmpx7ObQ1kRHtYd0R6JyHttIf5IEyze23qiabhCw+7R3GG6vXXAUIhfTX
Htp+VNOu1qEepRG2YJm3zlQO6B9ww/YTWvzAkjrQFn0iOjpE8NNYv90QDF/pjf1O2AJITPOrDY+l
rsZLOtcjxQBQNd43ke2XIF07zuj/eR5ZhDMPTnYbiRopIXaXXjTh5WWbw3Szfiqa+0eOHCM762NQ
la0XzEN2Ycb+8YDqElfZuM1NCHHvYtQp4npz3hPuzq29x1jDHyiu3+kYqi9Tdqe/f/3suaaCemAo
UXXKTDQBKKzj8Hv4E5KVnzbDbGeIh6l4FbczpGrJZSuBaDlTrVEc00Wcv16/irLFWdA+/jtK0YJ8
e16MqHGDktddCEKag+5tEhX0totpwSUXxxhTQiu//O6IQSkwtFP8K4XKQ7/4UunMMusKvqKcMj2z
dPQ2WvXY28778vphg0D3c3PSYEknuNf98xLPkF6SESH4vkHFBzf68qWqZRPnYBwQnir9hFVPF4Zz
czWpmmE+pj6CC98VS0s7ztQBrJ+B6duDm8H9pIL/Ukq/7g89nQNYP5AEjJXgT4UQUusi513p0WPe
G3Qw6IdOCz+HZ3+puBljHWkxO8ctJT0Mh2eO8Ba5lhG8McvhLmP993R2xPW4XjgWDIHaFuD+aGEF
hskPTl9sA/RDL0zW8bFdpkM6+mAKlp8MSgN2dIyD9kjMBuv4gN/HhOzEGGzoZckiu+muSn0t6ODj
p+4JauoTXz6BlXyv69qkKqqd7vPnTlr773Y4j1Iw8FBXB595HZOIPb4NgzwXVGHiQWKHr8uTf8YO
iUR+iTstmiwbqsqybrbNBQIo4lODSrUz0EV8kihNHJf4kudRRRea+mMi+sLrNvrhyYOYJT6o83CD
qt/0yAC3IoH2MBwU3lSnZb+GfxUFLUSpjkrcQ6frwH8xgZECuWALdY2aWG4Mb2AXFrV/MSYYavbM
CYdsnf5+Xfsa/gW8Al/zzb988NH50e+2Pnvni9zpV12/NjDBd3dxpz0AZWukERjtKjufebUo6qsh
RL//euNKO1Ga95PncDxVbni/C/GuNvljDLzpk4B/wXyjJWpWRvEcYhl8yIDVUppngzSrA81dNj1S
jdxmySgiKKjojC/fmMu2ccBF2HUY8a99zOZGoaWna3Lp4gtAPYuWtd5t+6+VIXuajH6+kD8dFMqe
o093oLMAyYMWO3CBj8WQDJoG+eDJBl18rXCfZdyvw/EdxflBJVAo+LK8an6DWp0Qx9jfGPGnL36L
P/OQJtWm2aBBzyCMUQ0x7ohw7iQWW0NCK99KvpR7UjgUHVtrtPed6Q2nNwk8hNm07RSNFhX2cS6g
5LuzvoNySH2oYl8FpO80r8e1IKBipayuXGbW/AvXxUZbCbAK/TazFpwnaPwdpBfz7hEpm/PNXY0K
roPv4Dvo+qCIcEc/dH+LFDToEcq0ire1x+BKxhTjLCXs79l7H+Vh8e9A9Wpo5CkfK+LB0aFahoda
ewSmEVFXxfcIsvbu3iKOLx92qVDLUHzZ1GkXF7+wM6xrm2aNCYvbBrpQ3XtEPNJI9wQhDwD97BHI
OJyfKUV3FjAEUG2wvZgPFf2SRNIMOof0CQfqn9I12K18q0f9gI7iO+vEkRwYsd3N3H+8unNgIXtW
69darDwlvj3Q95IkbvGQOJniM5WNN8noa8oLLaWm00G3n3bO4fp68yrSnuja7746ywhp8nRUelZl
pwFZRqJz4avu1UC8FWHEskgLnj8lfU5D7d0VFpJnDYnndaudIkvvZvMoaFLKCgVphYJ85q1CjFST
mz7hcJ4mjg8JV4zNbfkVdb0VsTLTnWDET843WT4B5LiRML4QjGGQrBvBUVNCNhukpQ2jbejfO+Za
s9w29MQ16O2MzGZKMGYvkED0UpqSbLAUuZhlx6OHcMbP/vvCY86XqPekdsMRdU5wuo/bTXx8CuPt
hMU1Cnn3QIPU9Tq1sjnN2X3UrhZEFl/ldYpuzhzTFk409BNvqnjbdCboPuQCuSQB7L64qkdc8qlj
IgCARSmjQlx9ay4OXBB1P1wdgnsogGbJB4TSoIWt8OEuuXvockCUGVcO3lZVQiXR9KNlI4lEgSR8
XsssENMP8tgc1sTUhO1qKFOmBmSW3kOqGLJdjOf3DqaihJDjBE10HV+eHV0VWllHtymTCqOhrp05
GvY5hAF6jU3yK2j2AgaHGajxeiYyMfJJhMo3nKTa87gDIlNW9t4xQjdpFIkX13EtOS4cjftX1qau
UTDhMT/4riRmaGYyjdDe573jQir3ZJHZb0SvQgoCiKfCBfMZ6m4elmEZBYRHs17HVDq4JtYnFJDF
+FclNjPoCqDMrZf+JXbydZ/08BHYPSyBuAg9Nv/37TPWFVWEFh+barcsL3o7kN/WTgkcukirvhY1
1qf/2M5Hb6Y44b/aOyzk6CEOtNe7aAVg8yKl+hGRFrLPBG+wIX5sjGH/oGdsKP0+oIcNUfhjPA2z
cuYTg5FWNKEWKKkB3tOTZqbElH5iqaF9X+o/7/w2P8b7PTXFjA3ZERgTnOvJpYV8tyXfcMvinlIg
mB1UufCbq5pugP4LNaekyG0zQiT6zIKA/5lCCbnPmyzXr6CB5MGVgLeYnV4l3PDXe6Bo8N+WZaVB
egA+3wmfkv47yJHe3c6o5ydBcsLBCRddl7kfuwjtEjbrQsfN+1DOjVs8T00fLFA3Bot5KhGnlh3B
ZCGAtgWv97MytTMufRonBTr5YscL2s6sbgBIr96UmaBpqLcEiveY2aEGXFIYtdvowDtsXV2m+6ir
GaCD2mZGEf313xGupXpy3mN7MyAnS2UGUA0WBsPe/nCIFJCg331Hlm+LyWoC8gDFNjynMFHIOyxo
vDUb2Lon4ZWulBNZAoBklUCguYA79jU9IGNQe4i+Zh/b3WfwGMJquB6wbHVOTUQf0cQKCU2TTGYM
CjZ70oQaFzMM2ckJZ0GJOm1CWxtmX5Xi5bJZpJ6353Zlh/072OnwAmNxjXlwHr05KrmPCGubgB7x
0OHaxTTdA9MoLUl+kIhO8YpKKhvi7W5Vppv2XoS7yB9Qb5XwD6K2goYPhcX3DubRE1c+/ccvPvfN
shMEVQxEiqEfeVk5u3VuWrO/sjGfpxq1y16K+zmNmW+/JQWTo5oHJep9YlN2XVVUiRWDFBJTLIUo
dnOZ7wLSFOT0Qy7zcPjH+lVY5JhWd0F6BeuHUlSAHUZBcUhEGFJcdPRXUXXTzhOo66gGkzqzkDZ5
6negaeu8NZFLa8dHYPVshDv+lUzTpuVNU3oa1wMWc7J2ZdWPenqTNo60Kt2zQflDU22hCZIRQb8X
I6CjCChDBPAFM+V5RlL2Emyz8tIp6aQ5sEK6jUZiEfMMjwz5J+CbE/P2E9qnJbqbg2KK6foHRl4S
9VNiHiM51zfYnkHeoTFDRpAn11dk9cqn2etcJXnov6iXL09WVxpQ91ttaTMX22eoK8k8NueiU2HY
UKfTMBBWVaHp1l+C5YP/dvMfla2k5Oq2zqkmBc/+ATobkwRo/f8OZwGQpDvU189lWU53Yre4o0NS
YQuGvx5X2ljkEzuk92mJhnr8BnD78YnFt7phWMJW8AoV9Q87gsjpQaQxGyi/spuY5yY+B5LEMlYl
NetkGz6DF/L4FAnlO/UXdGWdMJh3lAtAcyXdrQGAubsN7CvqMq/wq/MbT3XqvSORsHhM1ZNoOvgI
liB/CI+sg7ROGtezVIuq4PN/g240MD7V598/FKTp2Ik21MZf4B26X73ylP0z+43y7AitVDqSX1Oh
Ld5ZlXTBBtfCTQ9RgO+XZhTIHNk9q9jOyWIFDOxCxTWhTvP1xW4MOQ8aL8M6eoG85IEE46XT6gFu
UtssK+Rmeay22zyuNAxc9up0R2fzkEi32mkoRWZsge6GL8Z9ag/+Ervc5xGqLfYONgdY7KhJLASa
pjGpnws4X2VqchYx8wHasFF7g/KBNahxomJiMZFnVG9LiNxcjU/1EI9O+XQITXfYb/iiZh5ZY0Dh
p044I4e/9BNMNyUqMInDF8H5STGmxcLbsUpkG2cBB7/DHUKRzRjWFunrNulCdb4ZLDzeRRsGH8vU
lwoy7BdBjUNY9TB8/ogLA3sVuUwQGeUTAhHkNYY2UtaJpLMB8N95lT1s5N4cZnSDIZPTXFxUmRJe
1yOj+EbcvoLCudXwZDTgvU6M1wwEutrNA1Ge3cMexNo+SMsoCutPGaq9Arpl7uDGGQnRCGJC+LL7
AuWUoz5lVqF6yEXRr3Wh5sJXFM14is4prtzEljb2ECGF9YjqSDvznjFQTQNXgJgOt9OmPMLXMq2F
RJh8M0JZ1x2MDwyK0BUdNWqQGdBW5tF/FxebS+I438FUaEo2n6lxwIgh0uRRoOlnS+hlOhTVS1nB
MjovAB9qeLfa98Sjf/KxexathjXfHpB0jihQdYQNZ79iFr3KcMHvJXeCsbUpzHSGxp1wsaZ82KTw
sPcFlY8qz6b4LLPTgIpM+4GPXRQsghh3v/88qaY5sbFhwY9/ic3t2CvqdukRXpu2RGCIIjkRTK42
mbZMVbKdj5MZVL6yhFGPJcsKXKKGPWVhYPmnamE6KAyIs7c6Bg+8UsfybVFNJrPFKXKvWUg0eThR
Ego4PimG4QfOlR5Ios049poSWtzsQZrk+J8XaKBCu2eoDOFVQ3BDmPDoidLFKRyH2qsBC4MSSILa
EubmdjEwdjAQNAeXZ1sXO3CyMfNwxBZvAE4QHCzRNjIzPFEYAG40Qq3l9ZtvNQOdp8s0etbrwBzP
b8Fler3GS/Yiew+5MLvzA1c9a0+aJ0a9+2JVNX4vFQEe2DJpXfPKnqZwu58TJcItE9nm7qbg6qh1
Ana7nWiNmNgf0Yify+FH/ty6leOUEyd7Q/jJ+VFudiHOyxj6c/xGAGupH5RGb/AiL6lfWTwvK9w6
L9XfLWpv7VkfinD5a8IZtUpFSAk9AEcwNblI4JOPgua4ALF0UopbfzqSJiIdLjbhUFMm3n9vA5Ji
2UC6S3C2hWEJvekjowW7RkD/8jIYJNwGZO0tsSLVuKfE/dW4/PcQzErvEC+WOndr169ftQlbUG1X
yULSEBu6qaojZegKFN4v2JgPuK9WQzddzZ+sTEZr7ueALRu1fWJjoy7gSF+5JbufRbEkAYbHfgqA
SnI/hMbNMW6moAljc0iM+VGTQmGBn5HLBUA2dyGmZunB/k3y81SdrHlJ0RgPUxirUTAtxXdMUeSO
ENk5pkySUegbDmh998wWEVdgY0YeE8VI8ZiJToYrqdL3LFVjtwILlMqsFy75q+q1Z3nqStVK1Nn2
Kq9AQleZbN7xNUWgP4k3MIwyX5znsSWVepMEnBdUxhl1QFFt2KW8YPmKzcrZ2SCqggRogFxHdXyz
dY7w1vrFVTuhxXOuJS4grJb2Eq5qdkEY0pBGzsvh251HRofOcKoZJFBoU+XyH2DvuZ2RlazVGmR9
qOhhK37qaLLUGk6+UqA1rkH6NG7lWtjJDIGahuxnMJFsmGOMHsfprsHj7v/EfVViENecbM1uVj5r
54NiYsmhOqopB/R2DYwIcsV+IeQpfQkVOYJNrh0wj+wRcDKIbaTgedZx53n8e9X5Gl7aw5l1p+MB
soLjnzK8zVRWjPOHfTte9HDLG+e/osVGlO3I0+/x3ghKsyU/wPIxMNmiOu7tIGSUshaybzzvqY7l
9qELYKknhWrIdkmJzvQ2+0J3a91v46uoU2nJsshFR2tbsg6bJZPwM2NmL1hV8lAcmuiaAXHvKcJL
J0vib67CGSBpk1dWGf0F0GMO+DGD5Igh2xBWhWx7vMg+HrU+JfEoZBL11xaA8dxi6Cs0oFV2pQB4
3eDay+1a2TaGxtGZSJoomdy9CkmKsecZ13rfcNDa8jrZ1FWe8M/Tidrgshy8jEWbS9zNjgpJfx50
USJGSSHR0uMMeKNzM/ew+zcydPc4bXQATk2CRTOAcUw3P9Jx5vDTDONzCXFZfcPi3YJl31HB4Q+k
TA49Kz6+O2/gCg1dPNPtGWzBqD7vDUydvbWD/CS1Hl/wWPPLYeFsJcN+QRZKB1BaoK8iOYcwTNF0
GQHehvtbuYNlgoCsjkhg+2VygGkCcJf1obr1SEErqGjAQtiAAIQAtoiWZ8F88kiXnZ/pluf11Kxh
/F9n9e/CpUjiDsV+8Ek8OIUA+L2sucTQ6Q55qrunmRpU5AF0mGO4cXyMLm2m1W33os10fY2WyKNj
M7LKf1u78lTPVXD/3Qm0W3bVqaGpU5D9Q+t6qducngXJIbBUXPImVNF4HGdOzluUh9XtMgZdaE7l
VeW3Ve+QrDZo/IPw6YFCVqYgLAkOXDedQh1DovvKgrWgsgz/Ei2era7jyoyQZNCaDD2WYOKlM06Z
y6NqQQzQnki7CP3hojZvtn7PFw1GC8Zta9GjimBc1jjNqgTYadkL9kFWImkGLnku39q+1zv3xese
1c0xpBIf1kuE2LnQ2OYNqIIhPF0Ccz0NMmELhmbvy7BVkEBUj0g3fNTcNZRzTrKrn9qYwTYqjxXE
qDR9PIkCkHOwNNb0SDudHiYGJvo9uDnDjxAANVI9/OPxgRR2ZGQqioH94zjuhAU+zQ05O/EUOaTP
QozYchL+lcH0BQvOS0XasvEmW2OT7ZBCHIUHtfnIl61lDClQV9bodNL/5tPsF3IB4eJA26tD7qCM
P7xts9OEJjeTVeWrpS3yu6gITFsV3jnPqYOR7Rf6v51ZX7CNInSmnfKiSD5gKyjOF0iBHXts7tpG
BjlCcq86qEs0OQXy9EajheZAMw7opA1gnHU4uHr/YGbPSrPyue5UwMyoMYnOm2CE1iZfDEUtjujE
Jxp4MrrT+zegZkhKRSTVkyLmLtcSU+BB5pXyCp13Bq24wEqYt6CAoQhI41dxz4wv+n6hZD1v3lui
5Bx7j60sgZqCnBWW5kq7sXmazJVsquHMIHRrKpW63s6SGtPg6Pb9bfrV2xJhz5IgMsaPBFyIV8Zh
BRATwjCU3sGptwSdD07GBM68pojSQ3TSBeBtvNpcJnpQY2A/SO6YpkSWc0x3ofdTJLS10LIUlApJ
LrUiN68XQAUZvGHjMrJ5owIWPDDQjGcpiOQQ5mJxO1c4+DWD2f2zkwQuDHJgl13pxn3DpzkharLC
XAIpV3DvRjUS/L8QyWNgdj+BR3zGeuzw1O+K1TNJ7bHo58ieWVO7VyFhV/AqRPeS2PzRRKPcVtRQ
L9QnmjzpyCKPoPBXNn706w58aNT8PPmZAQwZZS5ziSxgZgaFB8tS0HYtQL+MdJtwXjjMZMuzJTPB
x6y40m5TbiOV4v2iHEB/dQi6ef3MUffi+LD//TQ4XG1rD76VBAu9BKFllvF9E5NFdXO8hwNfjvI4
oUCmaM4c25gjn+tc+Z/nk9hyhntLRMpLsGxVXQ2WyAT4MiLqGBYLNn6ilWCOJCoQgi599M8Far4k
y1zfQJ8qNcy5qXNWckIWahXzf4kVd5aazKt4Jagt+xWUcq2nnYtO0Mp7z6btuNWOUGUg+N5Sn9DO
Zjht4/QwTExoQQrfh12nS4flECADsgQQfOUREDhlmeaFXck3ay3hAnnRSKyZHyMIdkeHuBj6h7aH
zfTYApfduS+JgJSiU1dBN0Wtk8VwIx9u0HREYoKXHgM0EMzDKjm7KaDgTMi2AT5fJhXd7Kf157k7
x0UJsC2u1sp2MmdG/SlBffVxy0VNEoN16FVyL+300fDF/xPmMm/FqTWjKongOGd7SVkHySXX6Seh
kWV3/elvIrqrFVVWNdyTDhR2zT+Al07Pez4EEakgh7gVralcqFoq0W7xglMW4VY6Bo0rfCwuwEZ9
WaQe/wNu+kAVGbQkHihbT+S6BStHKtbzAPtN6RJN0TAFg2IKhZIoCQWVTnSGjlnqpOrQCzHRqujH
a424vINJYHAteXa9j9TNpw4i+4/n3yDsZL4XWOHIC7gCxbMCTLDAF9wdP+nXWCv/fCcW4mnJgflc
ZTtjv7+A5cK9FW9FeWceDZ1b8B2h33ZZyTmUSK7qWNHx9VP+F8adOE5nJBXgoYGfajmvxzS+ma6r
Ke/NIpt0QB2NqT0xxx8oG4Epc9QDGnyg5tYR/CHDkl/pmeDQUMXEGZOMhUZbzvjUxeKSuW57uCFe
miTsoeGR/zMNyLwkttkbpU6vuHEYjjnzNm/Ik/wARrFQC7McVRcQR8y+nTdH2apPaSWXy4gQtlrm
kjQv3wmnAWhChmacHqEC0BRRBQUOENicfKdGdO2neAdjVa3xustVyK9o/tWC8fEYVHnmY1Ny4T/+
OGB4YxbXSlGvODGdPPvyXoR8fmFrk4+T/P740XkPT6YCVgLQDWnqV1mSmasYsOAHar6Y5JD5VADr
VWIoNcvaa+btDgssZVLGOhKflptsDPtOet8PB4iQr6T773HajnqvtrJqLi/hrjeSG00ePkzACCZ8
ecwJ3BTY1U2RjOHhUZ+chFlen2SnOSvnwTikiFFe5Bw/DweNnKcbMidpWyWDquRSYxWwKRb7PnAy
CXqiJb0iW9GoIBX7Tzy1sZZjZL9Wz0tj/BYiCvpoJDxeYEo/eNuULNNGWIJZ0jAtfo/o2AxPis1u
BmCEI/icjVyWnPGocHqU+CcWn7ePePyfL6Nz3cY0GkxGqwLyUwgBPNdHk5KPeFrZbGxG1Pela2Na
sQci+LPqdUNKQECOC8zsXGlQoa0epIkAGrpVlwV+8L7KpBFqbOqWKyIbZdMWh64dC4Yo53UxK5bI
Xs62URpUi7QI5YqbcSlVX2uZNbyf3T3AXXW5Wv50FjRWYcE+HhWgEihgow2BIrnuKUEk1Luc+GbB
AHdAUkCqmuYNAgzYYta0ACX6WOClS/68+HjjOPLR5DnTQtRF6367Gf+DfNIBXeWjQHmHm33zDkX+
eHQIMXoRUD2nVzFKaG1XitONHNxBKoTMDosb33JQTLh9c0Ai0LVyysmY/y8LPLUcUkpRiVCFkjUL
/gWGSNc5BcvSi/MbKeevhQwBPs1pRRfUuEWmwXBkXLCpLjD5NnRAXt8b7Qx2UrUN5LMLJ4LHIj3Q
CuTSJ8Cg2+zYMN/iWPDY7eVw61UrGL6y0EXP+OuVc3RgBoxqem71L3fnp4hlAgDLScS9cW2Er25g
yao7ScHov+nnmgEpE6MVMeCHC10i/qbzEV6l2yLcLJdYWsHX8OaarpJfSQS4ZqckkPmh7h5qYLcB
3Iq+DcNZrEKhGEV/xJYqhxedqmjeZ5aJtaGWj9eJLdG+kONycWW1SGlE2rUkQOkNwVNK7v1ryP9T
JGXW5SHOYiq3eZZCruKMeggVBEBbGj9+57HGxKQgshYm/tr5q+9EZdDsw6+KCZZloyKR+to4Khnv
WkNVqun6yrKmBCerNIpz7wF1pcqy8ZVOM65FMRR0N/1dHeoRyvBZTAn+sUZLO+jJ+ln/lc8V7inJ
ApEc3aZA/YxzzUTIwd8vWVau+tAOr/hIR+6Ki0RSYqd+GYZdWVH9ZSJq7x2eHfTINqu6Gf4p+gjh
Qe5OM0HPf+H2XbXA7cWOKtC/NRrWtHksBYPQQNZfwK0Ihm7w7AofdiJkULU7C0pJ4X6D4WapgU55
m5nQDrfObZ/dsQnqlRyuq+B1PZzZPBqLxbfj4P56pao0ClRC3x6B7ShQggy6H88x+/9qIdZPZFMw
mXamtINm46MgkLHBAO8V2X4uFVjatZt2408NGcpWliaAXezUlmNNfp5EAf2hRnCzrb1d2fQOGyb9
+QfJZVbFv8L7K8D5bnwwJa7lzX8ZrV7OZiz0Q5o6V8MoPaOER1F9YnVzqve1gHQacME+FEd5fy8c
pbRr3g4shKa36lM/Ga9q7tWTqNmeiRPv4btDgam/MVwzNklX7ErvRaMDiC68X/KGEQzogbww7Okc
YND1PU3RWEVeeKgOq1xqTXzmgEIohZEjSHm+RPIYK+UWd6eVaxp4JUOm2Zh76pQ/sDueBuNDdx+K
cZRmQAJb0/cvvlXFGAtag8fNoHAPVYBSgItCYWk/y/jcwGcMH0L0Vtx8jILD0ww9n74yvVRemjKA
uUbqNIPw+v1cHYeJX8i7aIUrqSI9NVxhdhPaTD02SYQy8TFOcSLAYVoKRZfCxy3rB/dVZcsa4EnK
K1VVpgwjCJJIJBO5rcFgFIIOBsoKIEyq2u/3yf2VGn6+kEnQgLb5W36l1hDOor2lfywhICztRlKN
UB2TOYbkjsFpFwr1fRn0eTixzVS7WnJrq5C/1NwMWsvX1oe/MnCghE9/FDiq5o7/aGvtBNiNtb63
zQfvqGy6STbOTjnhE2iuzeQGujzdOVfVIHJfvF+vL1qejK7xJElpD9e/ZKR+lJZAZQYuauviU4wj
9RI7r9FysSQTJQqZ5GKuecayXuzSAUxrT9pV6erkDK+tBePTrtZ0lw7hX90f9OPykXxoiGk2a3lH
yPFcI3CjXbWWjtTJoOz6mXb8CEtb5flJI7AZ3WazJX205VRjlLriPclkWjRDfzv2vawIItL5jW0P
HC4xqvXFR4wzXjxpTF3JG5/1iNqQwMi/KM6wRuqfQAyufBavD5Va7ebDa8cIQydftqRMGKuj6e1P
9SyjRWwAzAS9ONF+/iM9Yp3mBBj42Bk6cRswo+o6l7xu8OP39GyGuevumoKwsMTWLM9JFsjhYclg
pXP6MtEGg6Hf4ipxDqcDuUV2LWZM3SX8nNugP83A+alor5kfDXS6SWRoHYecQ1akjef7/Z3JErEB
M3Ru2xsyLVtjQWdUBw3tUmuPn/pSYSIzwy1cTG3tclHgiQh7UlD3Qfw1UQPpreUBxetf5f9d0Jay
E0xE+zJxnJX5L03osIJV6VLuRAZMzlzQnvk3/HQ0QH6AbQ9bn1ReFBnsNx0felrXONLog+MBUqz8
cAXioZnNNoab0e8ZkWhSF/KL6yO8i7olxTH5TvqXIMjkoXNCxG77acQErQ3GWq7cq6essvcFFl6T
a/atNE3FLEkTPx4NpvE1McbiSyOVdPilL2ARNKMfWFfZ96epUsHXEN4gL2Jy5F7fWT5VgxJPEICs
ZfbZC4zaMKJMqbBUUibO0OS5Yt5m+9iQMy1lZ0BIMlWpWcKBiVt0GpFInsaZLtCRbFTwYDyBEX/F
5tS2xjTLvv8ss63KH8ctcdxAsGXZ4aR2HSWmYqOizqH6aT4ugbHYBde7XqwdjJoFBXkv+jwdXPIO
DlzY0Fu/LOjOidSFeqslZs1g9v4sCBWBll0ru5qjPmUQplCpgyFHClJXue1B11YWvfxJu6WqOAww
UnN/QKs6sGbwBH2Jaf1MosXc3rgdfO5/or/GHgDGq4aBtGc1tSpr3LLho3dxvcFemnHhxCOR7Vy+
nHFLqukIxlcG91xgThXGPRxpcYmV0AlM/b+OBL3VipLEB1/a3d86wgcvy1wdg2SWxwT9gmbYWsl7
4fkUCo0nB4lrxoxo6g/KD/j38jmFTLz5E3k08waWpckDnmGd+UZhqyWf3vufQwXXOa4VI3evQs9K
66CLQY+VRyVSXcDRBSgpFgx243hl3pp5o1Uj0bKOPdMmgk/cF/otPJSayaE7fY+9lm+dKh1xTQff
tdJQvOcb9UZd4XuIM/iZ5SLbO6kVoL3a/bAvPK9v4cdgnc/Q+4hGowDYxRwvh3lHzY3siyyF52/g
fZ4FJgO8t+QYTno1EXI32zWj56KQSJEZGyXVTY37c+6cf9E03rWdoGNGrLb5JjT9yDJIIZuM6PlL
TPEn++r0Q2XoTbEUcUWcczitG4I/vHWA3rtA3vwkTrKzxDHA2kjt14RAcbqT9+3aeVDGcKVFJZ98
b3uBpw4KJXVQODQkZYmVkCyC7LmF2NsEqSU8JEzhWmIOFZd7vZ2hIw6oZ+L6yhtsUbZ4UVqXjeiH
IdOak9tCLCX9dS+F8/pGkVr89D5Q9YHch+fo3KWW4JONDPZL14kpZHtc/+cUTDUzbSTEk+ZJnDug
GaTJDr3kiIZ33VVPYsYWBWUNz998HtPkU4qDCIja/PnLSBTC/8hQyH8hYMEqDy3gcPxiRCYNdtVR
kO3ENPYyWp4fylpSPWTgWOYzVRvP07sHTp+Ltdaq/Qw8s1o/BHJHckiN4B2s/ICZaOXne7fwYnjb
dV4rgHuYsrcXmUVmYj7Uv/VVlDhJ3V+QuDW764wkGC4HtPKb33LXJTIa7GeQnlJcBUem6mC6rN2R
HBgVZWBoM28aAwlCDpOp1EHPoNKMpJ6hT249KLipTPYoMxJL8SMfDpZG/lfbTTzBF3C2dzAu2dCk
Mj8ZSadTX54ofNYgU6iSg4xPcnbEWikcCD4FK0V3D88OeX7AafUa4tVFvfQ9jt8wzdbYuLnYrmXJ
nsDq49oIyR+OMhFWSUz1/tn/XcmF1Gg5QlGkl9yrd0E5RnoT/61T9VoHsLVV0RvgOWX8G7teX+C/
X28lIG3b7Vgr2eFEuL4iAnAJ/RERCIgqmZqpz/1aHTzHMChcTzcsAM3in8vA6f4zsANUoNm31V7G
id5BJi3joFgvIkG3E2x0Ji2Xn3EIXR0HzPPNJqOFt4FWiPCCwSqckhlZRIZxg0LSRXGjfMWwQIYF
PbC18xzARfpQrRQGa4K/JDqL/h4+K5TR9SKiRj55TL+UCR3n2dkilWLM7olNnNvD9rdNT5EXqsFN
ip8cW6yuZjZ3C7zpUrTPjhLLgvbaBztiuzuWMqq+vBzgMPZ9yp+OOgzYZiVvCqQkQSBzFBOAOPPN
RJnsrgq1bVIvM9ex24H92b5ZA7bLohUxG4Wy9s6UMfqFrJtejQ7OcSZ44FlnNs2lGptny9xFOoGu
yf0li52eJWsajapMgtvBqFFVTZy9cQhGgeQOGKaARboSC9ww2IV72156pELEKDHTo7zKTQQJkP3S
cO2wvW5lzIYuTWkQOt78ov8nTkocfnJX9FbB5E/8IJ5R/ukdopysmh3fK/1drzALfHgAYvuytpBF
tpHZOcQCD9cV6dN/hSna9yt9o71sCjg7j4A+xWdsrYeNThi1clxmpY2eX4Ad+mLykSNFePPODYa+
lOOwC4aoRQW8dhfKyRFbTYKXN1ZSfU1HJFxeqcwxbpFOQmYbmDXcZ2riBtp43/DI+/W5n12T0oMN
sRWZog17HxmlK8ao5M2dZwh+8PNrMoHVJb/1mAoh2nGP+uP2Vw8DbdkmbNCIyZ8Cce7AfpcuqBLA
s+iayy1OoWKtbPvXf76UwLxQ5vrwPC25gTHZjI4Sm/g9FVsnGmgktB0+dPIaWZatiBWLuvu6rnkD
XGJQakraKZ0Oc5Ld+EFp5ywCy9bZ4CttkAgO6HVtzSZ7fnWA8QNETJKYGB0WJCNO5AlXRvXrLGJf
s6btqrc0hc4wVn9eu3KVObbDxQfOzTxl68prwtQRpuIZ5xixry3hfIfMznoYO0l3D8W/VQgP/E3k
baoP+uqR75SqV13C0nfCPteVjG/PQAvQQaU9T7dV6ltAtUqUAh4Lva0KmxHSK7yq2KGJq3NBdOKT
2/eHABchqukn9tAWQZPkPvDxf6Xcu5k2CgPKUHJR5rKIq2BBq87Ok8AjUQnp4pM9zg03+M2Jksjh
erlIa03o47YBZpZOTCPLvxRtZnocm2l48XLIZqsyseSmlur70tRlPmG4vvCKfOqNFnN3TBqunfcl
rxSzFTsAlCCBqL+5VS+F4b+BPcSJ4zrsmcXDuiqY4eZxw8C4zuOgyey/xsGlGWZxTNNV95+b6T+T
6fqtmbjrx/xcPsP1GZPZn4aXongMJ/wgTKFJwmgNcsWa1mgRi2AGiPHwRasUJfgWCQv8cXMQhDKi
FmK/r6Vq55XOoE9uXLpFTvigZ6O+qn9s5p9jVZEFgbBl4yTo2p1W78Q7iKW6Qh/ewHInHDDYmZpL
VFEJsvd6/X1qRAehWIy2mfmgwDMmQPxN3v3Pxas/8tyDkNkAE64u9ZpWiWBQtjJGtm/UBpnJ/7JV
z4Tj0c3U9bQNJwp2G/cbVjZeISM9QoG5QokBj9+mJ/HiyTGOLHAQj/sk0WrYCElpLgNA3aakmlJ+
XIu24ZxP9UvETzwhpSN59iDqhLsTtIm9GtV8mel9EkwxhZOFaB2BlRjkYNkHjbbVAFamiG5yG3IR
oMcBMl9nQ2rYWidtC78a7Ry8V88/TyZqZobmkTDeZBFvLfN2k6achGNBmO2Umac9CMqbmLDOJXC1
JDOep2NbcUKaIbRE3cXMyA/ajt4jyTHQoIgtnq4ccibs2mu5kWYo58EAE7HiW+gsiZ4WMU7QI4Nw
pF9MUORyonH/tgT3p+cM2g4f4HyhYOCWZIfkpWDsBhjCgvbmNKPYNhufzb78kMiVNgCDxxkDD9RK
QTnfE1XWfNuwOHoKz7LmKQtb8B3QDy3dsqlTCWKDo1MfYKQ1NJWeqf2L6hjG812bps0tZ9H65B0I
zsIvwrCo2wtoJjmCUmagDr4b67xhz1SBohuIdWSa8bSaOhNPttMq6GLS2v2Y+lQ7ENm/wLyrhNrb
VnqQ5vmzkhL1yiiwDRDCGL347dZ+E8UzYBGLFYNNwefMwgPsyng+KDYiksMRniG+YB8yFw/gnpUQ
X55nojjRJJfyrtZNiaeFeLMz1G70Rk5cWL0twZhvKDhbWRHbcpPJ/CuC5u84pbQhN1+i2l+s02Fq
kUeEi5OheswT35jvlFeiGbiP6mwc3zih08Bpl8Sx6XYjRiA1YdZ4bdmM9dmmXzuRa/hml4ec+SUm
CLoXTqoJ1RhK4F9sjomGBpDsQR2/KuQAZJRoNAD97cKGeTaU4ZrUbKkw0S+G5OE9RD+rnN8kmOJG
eO++5G2sLLhZGEj8GPOEGVVEFyJtLB0AqWoXKeJ1+vEztPeubj4QI5vQae2mCOIaT4Etz6nRK4d6
YrPO8D3Ww3Z3SLuVXz5PpTUyyf/Z7/mDls3EKGpF7SvHOw19oFqpNP4uLlPOeIyqEHG9D5RbcTXT
nFVIxe6oOTX7deDdQvEHHmtfz7zlSAU66zzYuzAGaSfx9mk9i05gFXawlYwNEefQR68XC8jSVBEn
KybnVMUcjc2oUUiHa58bvvleadS0rxAD6faYJ2CgXZxrCaQuGs0wnMYAzeBxyBMISVV4scUjAcsl
zdfPzs2wY/yJI8XbVOdI+Dk/7UIwZNly8Uh1sTAjzMI6mCZIuXyuNhaUcbsv8Tue+xV4nm69Lg19
FPhh77Oa0ps4C6Cg3x9ZpDUSSNRsDcInstab4wGA5MT/5RsPQtMSMwIC1aU6Bt8HoQY+ndB/1uyG
JLtwpOcWwBidLjDyiKV3BI2o1Zb5eLEhyHHQjXcOKd6rZypp/E4uXcfvJqZEHEvuIE7FqhFCY8IE
G+HV6TYwJnuZ3NrUI4mgWfHDulEGxYDpoqM5y2h/uBLwydvYic299jObhvq6SbhLzV8JrJM3ZxgJ
DdlXzQLe8saiWGyNgp3rcyV/BvTs24zrev+HRrff8HBbx4+AlnH5WblUysF9a2+U7Ngq9O5mxDha
ttW0TeJdA4s6RNgK5RDrEak9pmkH0GnbKNUF0QkE+d2DTfcGu9P4qFsFFZ/VZd8S2Om3oxerXe4U
WwcjlwXxahz8uo812YjWgRbqsFVaTQA+SXOqoe7b1sMmvXpXxXQ9DzdkTGGMjXAi2y2AHrBE70EZ
vFvn702oYrY2T2d2TabZzIVrYFQIq3M8IOddDk0kHN+tpvNWjnPYvsqrNDQN2qMOC6kN8lrTu6Hd
8bWe1c7no9V6IS8U0oGsgdcDPgpLR3myqDmgziR/3wEyFyOagFhWapiQGVPZ3uD0m+DBYsyjbfbe
p4rGBH7zIF6JOXbxZLhZSPMSwPG5J9+Vn1HH9y2ueRh+9nnwf8VQPhdrEiPsW5cJTVA8RHsHZGHO
TmIMcxD7Q7DqrwV9+2Ma9LhP5M5rPwmhbB9EqoXZv5zUR4cwxML6+vPmzAU8gOKEDsuTTIOh5IXV
rEM2Hs4R+QBcXzY0OG7Ux1XOyuZsBiYcD4KeG4sWQDEuImpZe0bFt5V01vWIPHbNo2LdvBLGnjll
P/UyJhkPX2xmLr6rAj5qM8FmoDr5+048Xo1PTxvBPAxrjqvXpOCMnBKn7pIXccPqdJOpu5bgsPgL
mdewlJSRC89GHHylgmozjt7fEvNr6PeZeKjWv64xl/C0eT8ZoAJlqFXJfhly6vohkr/sMaKzCnhJ
XyyYSDwprg3aGBgFUyXJJJulxgdPRjHvdpdGK151Nur5tc/HJ1ZeOYnGkKuL1xjxBSmflu0jt2qh
wKulj9TGNF9LKK3M4kjyIN/oQOAswZPVNY1gQzEPIBGLkllArTIbd8PKPXEVI/dK7cLQQ9/MMxAb
QAmZ9qFmX4wb2Kog7Pjg6AYNd+W6g1U9z5Gldk+JzLiupfOCiC9iovg0acREDfBO/C1Y2x9Y+xbx
LO+D46p1WlN7NBw84MKkTw3G96pZWHEmBbiHuqqdmSwNeTGuZi0rRMtWNNrf17tZlBF1xWQ8YzjN
Oizm539j/duZ+U8o3n7jEOmY7Uec2WjvaKzizyvayXzfqgHiRPlzekZpmQmsl9aVTW+XJW/VXiOv
5MIQWtAOl4UBGifBiwVutmbx+C6dvHE/gyKwnoWBjei0orusoTF1rJpSPd6d7+rkHgdNPOXXUUbr
3UHYSo4LHNZ462xruuQJiX2BOvn0flifpybXTpIITwikEd3V4nuCSuWXjnYKFcOiNYWbnPyfDxdP
nivPn3XLMSXMveohZthpESM3gSXkcWyTYsuOzDbYgWRKcet00qftzKjKhlwYzC2XhdV1IODHZhAQ
OJt9qjk4t74wOUJ7LW4Z2eDAvzredhUuNbRh0jBBq4b/Bk36yszU05KvnhC0qyQ4cK42ZNIR9gmg
gchuL1Mzod3RyOeFR2HFrCFH552YfI456/OxW5tt6RwVcUAhA/iWNudoUiYbkGa05kurCp3ze64M
L4yBmCaNPLK55LtjnIz6dH9NGelZLqPajukC5OYfPY+vd5MSIdr2w0TObnFUbKWlsgt609xiEeC/
2V2LNxmOqyT7TGdBBIiFwblyRYWVb24K5EqpSoYdX8D82LCJflxmX/MvOmCyMjm47uzyPQW6ZKSs
wyYFyW80D9qWBOqxJQ3QYAZgxiR0XkZurH/KPo82I+MR2lPYSJM+pH8qLIE7Q1XHJZ3AiId6Zvm1
luZ8XdfIiY16zxrXRpcoN7LRHuMp7lFkYOPgCHfNj9xepiWsXBnGbtdxXXjySfGaMBL25awsG13p
kqjwKSGkZhKlU0VHqCtkY4yRV/XR8d0ZSGHjW7mORKrULjd7DhAIxAUVnBJJ3Yl8Tf7YR1r9Ec0h
PGC+pKJ+QhPCCC5eYy4aZmC7AflxDBqC0eneXgNE67cSEFPo7mXma0p+QwTXQIMmXYiZIsXV6JXR
fnq7gy802TWq+OpQI+EZ0aIVbEdr5j7VgCmBXj94yqskplXxUOwU3gte1KiDFvfHBTLkggjPz/yk
5kg3RzGi0RMZGUKtIEqrJeNfpfFzyoKY4QVvOUK1MJ1W+hIhWWzVjz0+xNVt8XZvjjd5KVgZfS8G
f2SnJU9Pz2FhmjhITyZGR7rfkQJYvmytYTgnXPDVx8Zp/u/boHLeHOBEaF1BsvJLpzbs5TEpjT68
NCpEfKSfE5qyfIv+ra/8iJaq7c/Tcwx9NXD/WM+Vf/m8wMdplrfedpgAh+KPXu4L6MA91D5kF3op
EEIxwIkDiTvj65iniwbUbvIpAtPmiysvpc/dXzB4t7C9Ku/dAYXhyKeS6PxNFUbZrB8Qfk81mJDz
oPQ3MTa7dSpjKEhMUC9eqNpcslS28HcocAqsIWx3r7YrsNv/gV4R3Iv4TTleZ9TAm4s7jWEu82Q/
FLrTO7otbSqgkX7NwHq5YoTUWPj/EMbvicZJYijUTUF/UzPJqT7O7dfC8xWnVFbwc48vqbtWYsZT
oMR2c+usBqT/NV7MHuYl1egkJUfQMwk7RqcYocvRRb7sbD3gNCSy9NY7MA+UblJChnwhxPcFzrBB
eyrq6XtnkL57oGppqpGAutblhAFkdhos1ewDK+Se/l8yQP7cfVvcwFqyREdwXlKUs/HZ5M0kiGqE
C02nm5Ctt3SavPCBB1vDBtmcARaQluJC+ccjK1WvC0/ru3GmZRyb+y3Y4yjbysWzc/GA49jJ921d
/6HeIJJOQ7GuxE2ehSmn0zsaReqSEZ0Z8hu6IHrM7c7imXSKwDF+2CV6WMaiVUvyOta+MO0fB3Og
cwNWhVfjq44Vu0TbYPTUdbipDBXlRSJ4jQaIdfe3XSHhah2VMbpmpOlQmJw3L8rIilbRTjPIeX37
FHu4H2+CJGmTZ55qIk5ip3pqWsHPHXmtrUDH+Whq+Gov9VfjwBBYQ1RvKhokf+IaCM1+KPq1ewKY
CClogVmhRADOAYmuhY9R6TT5QMW29sT8S6VXnX/sC3RgSv6hklrRx+V6QlCwmzLh/Q2p16KvX65l
b1RcaHH4uYSOuYnSvzukocA7R+sjqPDjCouyQpgNTNqPXD134vL0qRrKu2KKl5zcBjQuCmfzrKFz
f235uoM6O+9302mQWLdbgGdOppTZx+SF5hHfdE/jZwbFYiaL1jl0k/qN8G1uFfTpg8yJ9xlbTDiF
EaVQ19wGdvP/7x+QrNu3cOo1Z5VVZcMyWTcwICv9/vm7e1KLNmmPseHOw1MBsP9v1TcM2BVY+Ota
gTsU8d84d5aJFxER8Q8FztD+OMqus9VSaRXug3TqbcUKkOsAtJ+3oRZFwNEG13Qoj68Rg710BokJ
KzXrOiEhi1QBZ1TGC3ywlZZUCTyMqHLd6mV/1MBhrYSscOHEF7MRTK/5lu/j79hTlcL0zb8gaQ4n
dd+heex7pT6Rku2C7G7ybc5W0ze4QiLlf/APYkfvemQJ95PiX3ONM2zPI8jl2RKcOBjA1VL+foJA
3hK84XAx7ij5cyuSvhVGGdbg3yDhoZ7ourmNF/N/6Xu8y5LzJjG5OB8yzHygjTzPhkhFnXl79xRv
WP4f1aYgtB3HRYE7Mmtc7LhH8lFSHisZPkVYhhmdhjA49Q8reWAlZD97j+5uIqy6Cl8LQe8ZZk/A
uDhIOz0+Onl2ujVKkcCo+YHGkGdQtql7bI+BAqV4rTkgtbhq1zg5JUl5P8l+XnJZXPCyEWy3lmZ4
ZiqUS/6DekU77G7+mhoNKHi7l89BujbFrIxn+6aqT31csfX0AmWhlwMdEhz+DNh13uLFqmo9zMXU
Jaurm4iXx4aHgFPwbicAzTm3MmO39NVkyNFNDGjdUIXkogviwY6Yc0RE6MZvlKKRL+2h2KBIhFFg
ZtLAvhv+3hO7MVwkG5SZh9CTjfR+kZiZRJhpZ4EZtOhCy8ik3KLI+v7Dtmv1p2i5wYORpN7ht51l
BX/dD5jFat5mbSzPtNaNCnWVYTBm7GcspWQGSvOXRXM6KCW0iFVJ/WB6JasF2u7d3PW9zdjxNttz
PM0qX6Vx/p00Ea22L5V1eAHV/It0GHL+sBBUoMrqBLx6QGuWDga3pokTvbIi1lj9h5U/Aj3pKvrV
pr/3HlfCQNi6vA7kU1zlkuEDrUNDCfFZ3FyWblYRwT62QLVyYC/MMoXxkHLT82W+5sGhs9GDd6VL
eOJuMJqRHfuQSQKwAstiKN5NFcadWV3gcHK15dmaZJg128zQ1E6rPCEnuCmy4aL60F//JzYbeZ6+
R+SIfxIx5Eqg1UEA7T2ezbYnpdJUf5N3eWB9Bp/eLA2giZTQYXbo8wh4Mjklk5ICwSb6iA0B+vIn
6MJ8eVW2/YxSdnnhPc13ll2mmx+1mCRSTOG0Pi1He7TPfoQh0XG3eBnkYizhpZ5OxxpYD9ZihIOs
wFqwYvPPgrQY4zthLZ7rETZBUyAvgnvqg9Xv3P10EAo1UOctrVqSTCYF6WFLEbdQnt+yBKCIQLva
8AKlz8Ku2iNHb86bcN2V+Sbg24wYvUZbU9rIH/CmkJwm8J3eQsPiQjVFNTzI+1n77bFFCmMBjj7i
RhPaD88qhNOV+fgsSkRgFjxvcnGwj3n3cT691TwULHC1CZBcMcgy7sHmIQnP64JDz3HQSY5YxDEO
EPsetaMFoFTEXzoQwiCCgfAjOfykN3kCHwnnexBadYcd1hya0CvBaSGkJqZOg1traIejM8kgVzYE
cXqWT5oV/2ggS8/r7LDxw3QZIhhUAxNN4Kz7RUea6c62sRJHi6I0fabcIxOh0ozxlMn6FK3Jl7RP
OoaCvFjsbkFq4Z2pNedzmetwR72Fec7OL1aChajx2WOwr31iDfIffiQllWCqMvg0KKTv+AVWy/h/
P5HORfDDhMMk5AThNqST2CCmdQVHHkN+97LcENcWIPHDn4wzI+uy3akAKfoCTTD/MRoRmpqBk5Yn
K5buOzqL8tpkPGDQ1rpbRfSDUs92yMOcAiul+RBltZUp/h+o5X6L8581wffOjOJ6cqCG8ItGC1mx
YsOTZRUevvKMTOReo9aMgj7sGTpqNL6NrJy80gzRh214g++U5IMM0+OYxev+JXafdya74XrKVZJZ
Q/6QhTiFSEdJ0xtmuh7e4BbEZYROMLIol/11MoEJ1Gii9kgEHvXrPYwYKODzyl8xHVCGdPQVAyXS
cA3nTozAxg8WepQQykNKd+/72wYrcvHW1M1lxqVzW1yUfV9lmyKpCUMZ2+CJY01wNcfcgytayPnP
V+Cb/kjaMuFTQ5qednHPbsONC+INsmLq4NN8sCzw9u1+uNJ3pFB6abFUe9cIEQyHTwhf6l4muW6Z
Ba/V+LWm5PAD30jEqcJqbawSuGYCLZ3O7z9aNwSwgJ0sANAxdQhvBZOqP6kvKk6AhUg0n+nWTylJ
Rf9jMJOPDe2vL+fIkVSVXne3x5bK3nX8M3nBRQPmJxPKv+TqbC4vjALasms+v6EQvKJ1dkedarPV
Bs5LgVEePwngvwmxxf7CBYvho3upwTbtg0UAw5jQTT55s8DzzTyzOmwYHRvoIEhRbjfh7celDmq0
b6z/D2KWpwLS8YMKp9o37nzKac5/ZYXFLSm2qZX3mzJ52X92Mi0Og+SNyy535ZQ22Nlr9/HXPchQ
Rq2cluo/ZgKYFVwbWmzxKsZz7Y2aTwQksGWRrpLtRiMmxXjbcfReotC5+wisAro4KlZe8r4W4UpV
5AFZAu4akeV+UC1m1xO+QYN7nDUtqj8FxSgV6LK82H1txtBO3KA378K1GQJYpCXoAy67zhEWYj8t
LpG9KrVPaY5O6wZEA6rPBGy2mkDLr+F070tiICxXZYyS8Ko3loPYFnODh+7xQF4kwEVPHZ7SW1BB
mC215VmbgjuMXn5wiJAaXWcBfw+7JHFqtaXRReh6pYLuGUbabF4i7ieA4BqTMg7PBQzmJySktBdc
YPzWOSBGqAo9/gnC3hl+lzWji4HGynDM8rPMC0aE6CW+PCXpJ4qTtDz8GB8ufjJvIS7uKLSwi80I
cjjWx1WtcwpNgQJATtH8CPp6NWazkGQhYLqoGxeoaPdDrrSzbsXqI8qe1Bifv9mPbMqhdBUM+3/y
9crEBNouwyNnnfIFrQ1Ys5l2oozjQGIm5/9rYm3wEmfWJochQG7PnGlR2nu4LfF8jwYC5V5XAz81
tFQxCVc/PmdhFAhCc/KKBxHCJtyFnkYmj5U0sYRstRpoPZElWvVn/aAc2AHfqh4wN567AyP6bA9m
G2r4Z8NsuVtVSVDVUpbGsQthHz3OBJT18Y2fjuK7VXekjb1tC5ej1gxC2v2oZgG//10BLg9NzRQL
tKKuOtzU9vWKYQE1RcQ/rwiIdaaRYM09vCJGu3Gg+uUs+OFzytFzcwahiKCBvJyMXXRIf966dMZ6
LMXbL48Z72KWo5+zMgKGmN80+FXfZQ7CCc1WVTpnxFEA4jqd9/KYoveQ8Bqv13cfCtdgpLi6PUYr
lAsLxOhfTEaeLMc3rEYO8z3wQCd1giWUjqAe2gfL5sIvMlzxsgjo/sXdvrmimEnBJr28GwtYEVL5
hRoV5q9uB9dRfEovjA01f8pkTSCdT+Lzm9hJ4rZsoL+HwqZcbL3Y2118oYtg3F1WY+7hENh42S18
CyLTKMDZyzeOa215dGFYSAH1b9nfMJ5iwOGFDCnhIcp6ioMxoXTGJD2pHmJ6rpW9qiGElVuONfnc
HPTdYbWsv5AdoVLPkrwlkozqxfvmxa4ZEorhtTVdwLtScWujeAcgGvFgXWn1Uadn3aE6ukv2g/dC
M5mCIRAgnJMS0wpNl56Zd3WQQvx88j+4fLxKF+5SO+043jhu2dJjlU12oLwrSEc5NkIFHjSuvhlZ
Qp9oRbaVKiuNGhCk7/0ib3n/Wp+xsqWgHlRnjMenL6vNp0loDHjPPfTebm84816Wr57G2NWUUWP1
n9kr4CB46iINXPBr+IBoeLnHjsdAUWaF/K60yehvCNnNtPqm6rXX1KGTt2bsp7uHu+qWgdpfp3Ko
UzYQsZ6enDmA+Pi99uWk7RFB8sVHom5d/S65FCXZay3O5xXj4oiuLVhj5GoBzJEIY0olGbkIoaTP
l4jqnG5560Z/bspsf7Y6ux8wRYsr6orxh1zlXmVPXJr6JVuN/xJYS75R15iL7kZTYW7Gomghgun8
CjlxfsXPFJstturh+9SDdP9Iqr/FZ24hK2Ymr6gkAXXRyoC48UGc6lenB+EgJ3YB2IuhJsG3FxZk
nYdiRvhVOmt8ECeXQjTVqsEdrSL7mMsYcgFWo1C4mcZGR1n6UlM5oJLn1vyVu23zRTL68qqVEzVu
qNn7Qvb/QBVbggoz14+cHCPV5FoFh8hs/AgfDHHc0PcaGt4fpvBkP2XxJxbTbND8GvlxSLXvp7LH
RwA/BBKG6n9LhJ/sqFUpp8QX18O9+fxBMVAZSQ0WBH8Qs7fw4nSzY+epQywT02AJ1YjXUEpntisi
yHXlWq5hJJV38pASNZP3WaiDQj/Jc+zYbSsLUb1Vb8NukElB62ns9QCSdcqbmyeJIi/hbHfL5Vk/
grkvvJao2X9NN+MHFG/TH3mf/QyyAiTdhrupaDh0DA7lZQm82snVTQxIRf8MjFyinITbmzozArRi
VHvWM7VEPWxAc0l9LCNA67wH1LbZRqC7cvrgpS5nGIBFG/4cHMcFNJWNiB8Iszen8rc6xadKHJfl
VjNXwg5eZJBlpXna5l9wwpCt4OH5hf2W/eMoGV4wU5qFAUxtuOFCXV/1OOQ4yJNoHK48RoSzDS4W
BXPicH+kRYSVwDVY6Qf874kV5xNDgPvEMCuAutOz02Ess6NqVa/YMW3uKidyHltq6ARzIbfkaojb
3KtCy+HMM9VGKoM5a/q0Q9d6jjhgdm/dgx/OuGw6kxeElyxb7c4LplyPZaXsNirA9rOYc2mtY5aT
YKcFd3inP4u3FOvB4bLXCXCSdYR8Ys2GEPSuUp4JCvdX1Y0fqxatEbd07HJ3p7qy0BppJtZqOdk5
yeDZc/WyPb0mECylI5r5TZMyHEfI0l0mGV/Eh1VjdPmxcyE1sahVg0DoniEwFp2OHFS5R4XsP7DC
U1XdJqovLdLwOb+8gCizib/QVk8LNBzYL3FJxz+OnlS39zFfrfR5Xmz0xUlieRh5ZgCfq5hITIdo
du4dy8MNUwDoJEdNdScYYrehqHKdvkP0tqdG1QHaweMbNC2lCliqE39xU8MhLEys6Rz9jc5azPuI
fsZMp3G7lUFcjD0/XI+Rg+tW0H2nWN3hy2a3bbDC9U4kpddF4us7Knt9ugkQIRBpVhDdIEVZVxC1
OFvUniTUfL0h2+xL+Pr+Wf3IegQAJ6lI2QiQfCQkE6KFCMdr29GS6Rt7Kwr+dIqNAb/kP2bjD+ar
ec/Roa/j30tQSFU03eEWSTPn2BeVqO+TUjnsaerp6ibDEzxwuOv4MwWMgtcTJBANavVH1USIVAak
mOoE/Nw72gzv5+Oex5kongmj/5twPZnQK9zv84DRrmBTUc737CUND98kN+i0l/SWRilTHnug81Dc
jzn+qcr3Q+AK7S5zF22laJ2OeD56m10Wqx3PpYKhrtUBeIgxWIOzmdmJaqRelVve69BWBQUhWc/y
wDIMO8HDUUsw3JvBDAMUcibj75F3tqn382NwseUD2p/mnhShnkx8ZDxrU8W7NyW6P9w/CqXiXWJa
8BS+YFmdifAPGtz7Ug8oW5uFWyhbHe3EvfS1Sksg3bsPoj8FyAcXE7N71PMc0E8nxBAeUDLFUgTM
SsBQsv09QJlshSDMxxqAImHgcFQYGQRTKv7lmwYpAGFCTyiALF5mH+BPuYMgMRmnmozzQYsP1Rp/
EBYunUz33KlISvU/VJ1f9DLnklz5r5aG9WuHUQjIMKXrSJu44gNESuKkiGlkydR+y04LVO7Dslqg
GbY2wkiNqCMxi1I74mKZ62jBG+K6bpuHWBBbDvUnDkEcd9eeo7sgexrF6u/2JAAIUQbIwN09NPik
RCFaOqNEJi7Up0ehugJD7yVd69pqlFMOrXLjXE+9+bnMuqmC2hHYnYMMGpDQGx+5mxH1yhiRw7Wv
FXGrPc8I54bEGYHsvir0QU5//t5rvv9JZHIXkMlfKkDruSAXKA4RNY7sRwha8C0jDo4a326v/vht
tt4cYdvrN8eR4gcCL9NHy5gL98esFxUV3zEP9RFBAlqdm6ibFoomhmCT4y33oN/G5+L05h1Yjs72
Zro2e+1rxwG6BMNu1cO1eVeAZ/kRZUBJRpDOPPLsPJS6vXrQUC5Tv/48HBRVb9sQA2ejOpcWfRv5
1RPraB63FabQdB4wESR14wFuw8pz/Z6z0AzKo5zGps48a5Lnc2Wee0xfiKykamJQDhexsvc+lTv2
mum6NAbHFBavfIdTSxOIRx/hKNe1lbgUOfCMSxSEW1FJGyHi5R0Llb+u96iqfwTCUPURE4j8eN8j
3hEfS99unmpl/3DtISQq9vw+5DzhEjFrRZn/K9qtdEkeALtWgIXgyir/LHPG5ru71VBrNp547buq
TVwUFWZy82CK64sMSkUhzgYhFPX5Nk5KTJMQtqSPgm86A10c7+h5a7wL73E3rHIaN7pLNumENwus
me3kPFY9iktz384qHlUX4WQ1/fSSrPG5Tu7t06ZcO1C17cxQzEo5HwW0ksbeOhdVrVWrgzdcrxCw
svdJTccHKwBIa7anpnRjOdXuv4qjlMKR6R9BsVMGgd6aM+EuOhbgYLo3FhZ30o3Fm8FX2mXShYB1
iCj/fvmbkkX7UfPGnbnmK2CkIsIayoEy0W5eA0BXv0LePcbzpUJsKoHzGEKwwdHVPuV/c4vRcvP6
RWssAMrbgoIAmrasWtOkFjbD5sEAA7nMYvO3z6nAGSC79/xVkFZSvnLaRUMasR7XioIfZxXZVeiF
nc9Ron/ugl010mdQrLr+3QXk1CuT32G+Ks36jzFzsQvb6MhHUP2wivI6qzeAzPS3QGH8L4lka/j4
TY91embXIg2i4m9ne45hgPQMI9PxDUyechVE9sbgfrSoWtwvTSb9t9XhxmxfMbecEfuB2uKyfg+J
MftiQq8sMyX+TZG2lQOWuWqk7T/+7jqqNm/vaKmZoARg4RBc6UYlkRVWKAQzjv3DCFsDANMIAfmd
2JaXcgb8YTcUtGQjNhw8gTgHsv3uCmP+3HuQ8/h1x6VxkxcY1Gk8M8tqUg9T8BKe/6Wl8npJVbJf
3swktbxGbSajLzht2yo+N/+EcvlEjcAXS5qNRAvleA0OYc2XvsFJYa+z6pweRrwySBpy/tsPSFD9
9aA+97C1tY8X9vDycWnGZ6n1neELYe+7roQERqrW4xbFD96t29DBoBACsX+BqMlSUSqJgajGSLLA
ZGdxg/1xIzft07tcBmxgUFtqw5Nw3m8BXsLUSgvgCOIqAk4oQudNndJmKnyOjd+2XaCLbSGpo9LC
HPKm2Cpxn8xEsoSEfZ5Es3Fdf0t221CzoyzU1r9EQvu1v0vZ+HyXU9f4ifNEvoVE7Vy1aZZ4cg27
A2tJUEVrHPAbQXOK0Y1U49vRjvYGu9M3KfNrSneV8vzyHIorEu9HOQqbKwyGSXHvsDAihPL4rzbc
o8uatViym8NE/2fVHQ8vaARskYdAhe4qWO1QaVSNZi3KWXjdQNoeLrArh0Y3EbwvJDKHV+YDk5yM
MQLjVrpNbzqFdgLOZo1cH0rbPg2O/FKqtQgipDRzpo3ofqTW564Eqo4xsGrIzE9L0c9EgtWwFdUb
hll1EEpl3NQrWKQ9VewupIHjn2WT+4bz7s9nfh6BTqs8khFkXZdvzO8Dfj7A+emWYPQvWUBpQeKR
X198Mzvc/4vwLMp2TO0TecOx5w3+n/yUorH0jkIFW26L8Ne4DXQQF0FVF8gDsNKQxBOA5L+65I+I
aOXwqhyx5Q1he/Iy/DY8aH9IV2hpn5nAgBCafyNifW5XQELhIJb3AVmbnZcfwXYCHC4w9dVveBeT
/nZRdTIllCKAekYEM97EhAW/wocxs/E65PCHthR87eTCUdYHX1Af2UBiutUGC21pIZV4DM/Jl0yT
GEEmeaVyO6/U8BGS3hE4V3l3SBPuJnRzkbKEnV6vsOgAZ1dihZAFyWdam/PKDVabojxNKRQ/sOeL
Ilp58wejf65FuBgNhs4e42jaT4NceUa/syW/xVf7XKVi7ab0JXbfX72ILGIV5x3RFisaWnKarcqq
CGTPrarUbOWw4ZpxUyq9g/TWg1GeTd2zEoNprJRmXP4e14+3KcOzx6niexpJRSn0g1LT9GatziXQ
z1q8YQK8Ov0NAncSQ2LFTmm635N6yPESd09gVtzIApNVPjcs7Vr2i2Hc9ligaJBdE8SFko91+xwa
CkZQ9Th+pkZixuARD5S5GemkqDaQNgn6WFgk1tOfCtpuGJmFfPMS3JaqkcBzU/wJwfpyJtK1E+se
SpPFtuYZKLiURiFGySlHcOpAVudsYKVgxaChIyiq+uSfNv8SOE03pIgngcLx7DY4O0nDI3uDOCsT
AX5jUPi7dx2JZD1dhEalK65xC/JvBY0bNi2o4p+NDAY0O8MlJKpRzUp1NuGsepSMd1AXNVabqS6S
JFngbOyve44ZOes12LfJK6z/t39JVBZ28YHO37LdGt0HbbHiZHI+JP5TSOuMkyb9FbsSEHRujUE0
caHdyhPwctb8H/aTWa+FtjvxtEfX/7t8nExLRxK8W32+tFy3T96tEw87Objz5ntRrzSzCyqGWXFB
roetwOOOtNx2QBG58u5yrDVR3G8pHQ9+i8vtUuQ4QBEOyNlAj0BbgJZy+wNgviaRAzLIKQVzpkcD
Gu9QRndm1LP0gm4Y09Xaamg0UZLhkqBlSEdUKbjK+V5P1FLjEc4dh7hMJif1aSvk0R54pnHAvqjL
q/203AhQ40AqSRVrXLZyXGAXaQnZRLXueIz57wejjUBIneF3ituZesB56SrkembMb3kiAuMa5kBW
O6rRbvzP1kfojzr8ENdVlI2l9DUVkpkBVK5WPXxyxXI5Thew9S0PK0+uRtFYNqTCrDz0Ad8t+7A+
w/mR7Un0ZN8ZnsphaJWj8YIpYSXJ2i8Qd1t7yUGJKYqBJnd3zS6Hd3lit2EzVt6eoQRSnvDH2YzN
FN5VYOLNZh9NACaMoaFobgAZ/utsK89MK3e5AHkscqJSWu/WlHfGhHukexq4It1nZDzFtBBNm302
IWrJ0DFuwm/lPRkwktIzaQVSG+gdKh7th6Xtpb8lWtzJvvgcIAVWSV6nQlkSn7RiihERtXeZQA+c
/IXgBiphqKacnlMNTzU3NKjunBOeQl8=
`protect end_protected

