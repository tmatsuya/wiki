`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRCLQRmwIq9S1sjnqb2dDsAHYQHteDLgSVeOx+BLan4kFwY5X2+XCUd0G0H9/m2ccBwq1pqNRWaZ
9IomsWIFtg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RxNz/7Gnpv2owxq8+C3pRJfX8uM1tDKu1KvIBqpvYXC7roMAVFi5BYaZpiDrymsc9G3SyAtxwzn4
vLl7iZChSWBEL4oRHk/HbtKJg/PZm2dcNyr/jWGYVPDbzoCHun4PVuDhTq4XIMOW3eRsTk8Vq5hy
pY8otS49f4Mj1yLkRuE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RrOHV2SXQfHIEUYx8qXVFwaA4hVb0Uq/SWhq7Tkqd3fAXagRzXRPs1aO4zNtyNl5gWjIMJoWnSYE
J51/R7RLafSJb6MBhy6u5c6FXNGKNotR3sgYpK4xnmo8MaP4Xnr7saD/giBFcbCIRb997V5P8YZ1
lJD1c/sDYWyfNuLJvRnHdHw0mUrnD4UH9Dlc/FMGckLyzkofzvAbdWelZ8OPIq9ipS4btylXWUB8
z2Z8Xc6c0OSiEKr7izKSYSCHYIO8HfXgVqlvbmKyzVN7eGfNoDDg4+uSQy3B+nu9JqpA23ShBpaD
mPo8sOE5mFQ4EUGbUxDzPKkxy8L18h4zCOu2aA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kXHIDe097KztJ3RVOq2N1x2WSLnzzDhnsrgFk/EahaCQvGWTsKMc3mDb4abYu3STpcFKkv+8RWiO
tesjzu+d3dWo/LYjffEstEmznkK/eXR3q0eJOH77/lU4lyo0J5E5ragEd2RHp4FTo1RclKZhEeQk
xnkbdQTd24SoOKFdr88=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kl7O+LtL/KzLDsdRO4doezt5EOgpfvNz8KH91C8uViP0CNKDaV/qneUBiMkdYR4nU8qZeX8o3cp4
pucrnLNLW79bpBO6q4FQHbR6ptG7Codys9XSzp8HHqzIcZRXqnqSPAoPOiLqtum5C366YBYceVfI
OSRnXuoFtUXW37bUiwJFjydi1i+C/nbUmMEhuwdUrFyQ9SeIF+Q+4lIlLPyRnFw1y4qGhCyPBQja
P+AeTCeinFmD64vmg75/Ds67MC1X28mu/XeeSoVLVbmwQ28QYUlxrTQ2azUUSlgbbdKd/Lpdvorb
9r2B4xeINPmv9qYKbZTvaBHXyKBN2qs/YDJj3A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56544)
`protect data_block
1SL5XX1hTt0ci4Uvp/HXGNzzIXOiplPvx60Mt+EbqRpghmiJWKuM1KKQm/x3/CZiod7yGGebhdIX
B85XZGV7zdDVAR1pdiTcPr6P2szLcEY02mpAlBwgAy5f45xpX/5EPOs1KxmFHXtxR3/w+oYYurmz
GxZktdUsEz01n9PX6rEMX8BD3n35Fd7NuQ9NTrKOBTolWP7PFXJt0j8jIakQNtwIlHKv2xXNX7XZ
uDyF9ZoI0T67kBZDFlHuPcd3mspC2/s3z+T7DJfXeo4MdbBBLoyLxoYLuD3xhQYORvcOk4+kWRUy
h44RHFFXutRYET0CSLKSUsS4b9g9k8GN7/h4SJxIrj37fjXso+5/ra+hHsQfMJ/DnYl3/bYGYSxg
31XkiQscJfeZKqFmjzqOw0Iutjd138PdTLXJXJnLkYr/vGh9XVAGp9fUnDPR/h8XL3yVGfYWz/hb
++ovF9KdHEUeXJAF+ReQNGSiiMz7BRbSaOVR/X+paJ5n2S0SZuxOScMuJgSU5KojNWqtDmlfYIUa
QF2ODVwc1WzQsoSUx1g2T3E9vF5PrWggHTO2mA1AWdGsdIgrAIQ2gt11jDnfIiaHss+lZp9ysLgh
mMYqs1O6oC68ht7clTWRIR3cSLNv3TQnxnB+YQOmxuCphdXAwT4i6+F1dNqFS+yCe/IDnrmpw6zS
ndutL2+/sdxfvIYwvloyULP7OKEkQ1MXck+BWmQ4CpGDW4PXV+y4dfIQYZWV7TyewQAh+B7dA5QO
8W95OAZ17kXypBeJvQGyQHebHv84zv6Vxom+v8Ao29/4Mff39hXT2gG+B2b6RaoJHgDzy7UMtKRc
fIqp5dkddkf0lIe4OhNCsZfYostHI41R9tBmN77XRN5mqYe9YXf5wuS+cT+QiOOolHTVB8mF1RaS
Uz+zSejnNhdnRVWlyyk54wp8mDba1BEIXjBP1lwHKJWAyISiltXGvltx4Z8IG+eaNuqgNjlib7tl
uTkZvycwrX1zeH3jhtKqBMBRgjJASNa+0oS/Yztl++AFsiHPcys5/0+beP/2nSXq6wMvY5Bh4XGw
8qx6ZisnX+a5dSeUWfSbWb8CWlxJp87tLLkDwydLfzmsu5HtXrZXmDj1BZnGAWkmIRssCIdghOYE
dZnyvN1L3Iddye23Xh1LkgX+AzfOnpzIRZrTjTb9F9V3PBHjWfD+htLMXFf1uBlc4XErm9ZcZp1I
QYQKPal5mJZTy1vcpNEY6ZF+5UQiERKB5o0MdpFpFvDR54fHMvfjKLObatCOEZTDnp8sq2CIqgMf
/s0K/vAX79OiNeCX0VX6De40xwC7sHuzYAkfSzz46w+O9pC/DXtB+hA+kSFTTYMOUvDEjT7JoLgE
MFqSf45LDXcb20k7X4OapO8srNN88KCbN8umB7xm/Vhvd7dSDJ2thA4RyzThUS1R2snCGTZzPFTP
USYBy3dVPohFwA+4XyHWqBKA36Cf1gopa4VaKaLKU83ptJN4AH3tuYdxQd6C90TwYnF0v/tkb0FM
VAmgG4WW6n8I8RtnFeKsn/LbZFpzFge8K80/GPJdHA6rNbTO32ADy5PdT0YpDmKvczLYlkMlvf4n
d8jVIQnOzH3CA6/i2AH5c5AZNoFhTQ1Wli6z4dN9/CrQkc9Gn1RE8+tA5Dy2x2pSBJGpu4YXWRyM
iXj59P5UQEqGpRW8duHm4on/mHqXUVMBIYptBD/Vfc2/G/W8HN5lhp8ESbHsck1a9R91cSuKRf4C
BjUwdxG+71nDyNSYmMf0o2NPLlx7k5yoU38FgfU7Bh4Y5IB541L0UD09ZiG09dKf7EWZF70rsqNI
oi+u0ZYiNmotcoN1SywSPPt62Egw4C4yHOi/a+qh5ArTcJ+JEYAUsEZxC/zObcOlWHrTH47mVyjm
Zfnb/cY3sOCHQapujuUanKyRUuerQTYlkHCN4WbW19cYb9xKifkZNEpBSD6356cXks1ohy6QBiqu
uIdRyhDWAV1nFxzwcDT3Tx9HB/Deuq7sRuLjAVOFScxyio1K1j1GZfhC9QAmPWWXP2DgTWYopMuw
YMJMMWKVr2FT4yLsJmIfKUxYcHk23mRsBrC0wi4Gr/by7hKo4q20BfkLHiI2mo0HZAj8S99XEt2M
lyJMy/JkM2mmvcLfKYq+CumUGaEWVeejnuxcXE6fbuppEqARXHCRRDq2uWU3wNEYM8HguswQQbr7
iP+hYFXHmsqSQksRdi/epcjimkF1ofikvgC/m4fowDrUX2DcUUnIpHQ4/VZWuY8Wu3H/GUU3bcOw
goY849oDdiONCFmCBY9ZvU71CjWLzsxY0J8sdkQU9fxAzmBtgqBzFD4R7cx08xXGR7jzPfw/kXuf
7gRYoZSLtW7K14muGftZY32G6lLy4xa1fglYK5/JZlEkjjKG2Y7w0WADS6+N2+uNHSji7TZLZVj2
ycBSuxnffmMmyAqi+xybZG62gRYaWz1LRxSxL6ValFACIMjFkK43qSYg1kumqnMKigb+Ari9e+n3
kpyexRss9EPCPvacnLJkMBDId1dLpWsa/oSWp4tGuZL7TIXJBfSXYZHUmayrQFdzXVqiid7N9Koq
+9qTdWZHv04gMzi3hBmCTh6njQNVKfMWdVDAy/g2x2+57eRyKyxWlqyYPzXZlcKaWglwuH8xrNsk
sb8iW2Rk/O2OLw0bLP/SgD8sran1iwFGOLKCSkJb4HgsrOkKYk/MqeL6ASPpxqAMbCgETt7x7QDS
Pa3JS3XD/0m7rVqFiqWoc4Glgnt2jkf7SL2XoRnMdyEEYdhyTcB/SJJUm+UHXfe3AcmALCS19oY7
boYZ1hOHfvCaApnmPPButoFHK/Fs0A7JFBuvaaR+1P7vH8yljMtCOPvhshKzUbZNfbZelxnuZvGV
rqPVhrp9EW52K2Nlafo7obxN9l/6RZLKhQuU956ZmVNNH0xn30xsL4+/UwLmBX84MpxdUqLK3iKn
BlVc5FWVZ+uJD0dZDcdHGs9Gi4Uf91X+nPNTBhwh0mJORxREy8oNUWrmw+9223PpdW0vlbx/ej76
TKBKwHCd9O47gTKqjfX0wYAOJjSJUlW6WYXFBJEeF0U4HzZRyH6xqrSaPOMzghh3JPA5uVfIhiug
ycmP11HOI8mQppYejM9vHXQCi4lhVtz8fEL+uH7RG051n2+Dpz3ZcRxTVPt39aDu9L/s+3xTRQ6r
RqCkDo3ZNvEEeKmp6XH68OmFrGCQZQa/3H2mex4ZA5Pg3vNWQEC2kG2gZe86pBY+jkCX0cgZZ9iC
d+Jg64lkgroN2Tss8NtmWjBQsG6zs6cqzCO3jalNRC9w086hjG2RgcjmgnLAZOtS3yGgEaT502qW
1Adl2pVPeVlfqPnpvC5NO93Wi+TzRMf8X/wqDYVdqFt+bkRPq1QvpvdZ9WKRVmWL+LHAbvCfPEbb
itIE3Z8FziqTabwcPej+poSy2yHeEpGpRoYvQ59GIPM7SzoPXePn7WecHmnktn4r+AmMw34ZqOoj
FmgkNCaW8fk+/gfNhiKEFo2u+d4tBt2jE0uu8rSTAZQ3JJFKJWUYQm4tGDbl4uF2w6C1MH7dfLbR
Np1xnzXw25MgZESezFjSsYhIvIOUyXVUN/zZtQSfDudp5ihkQUs6+/9jkY0WgrvUy9hYrP8SuLcU
7LlcQvQuy9iIxg8J04FCCNLt1Fm9nyhZ7Iwquf2lC8ZyeBw7kUZfpAm0/ZkrXoK+4itu8IyFrF/I
P7iarM/oWXH10Er1CIClJ/WdMHsy6zCpIqss3qtQCgaPNorEHzs6ds30NUN/VklmMC6h5eKe+f3T
dV+Iy2lCkSZlhY3YL7Q2VwkfNmMw0tbTdHcYtB0DzhBNY9IKZoPqThWUa8UXpFGsp6nqdTXTTp0V
/PCCrAs5xcCOrzx3kvakcdNMP13BvV+wGPjgS0RBkYSMAk686MHEhg2h12K68TguTkmb6Xmxpnz1
tKZT/qey0qogUd4n8GIdOI+uCScXoev/lV2zoca1VQn4i+WtjChNeuVMa0d4UbmnMSfXGgHiG6BS
jdxdzEJbVR5T0ab7TOu40oB18W2ApjdyamSO8gvvXU8wPuM6sOvtxV7IsuuIemXsI+ANQcycyqTR
lCfsiApcovg6mM7D5A3S9ZtytK32zUKjAzLfEPjL5iYAHZh2x9TPXHgCAzCONRXEzr4ypQn30ZJx
XyKjbHQCzHYP/si/gW4tfZ9xZ59StbDFyHwmQZBY1wXLA6fCxKNuf4vP5XpyTbg1vlxE9rVjooMi
rdBQJmHhdwwSp2Vm1GlWSxc8oJBOFV06RRmf5EsivjGI7vwAWFUrWr79gZL+24Jck4YZOx0/7CC+
q6D7kxJICfDPJjFHK4LOyUDae1HqgmoLkaR5UXZYw25O6Wy9QnHaaZ+FioIoEwMFhHTxmsWZpGyZ
4L1a7k955TZMEnwrrB4y8c6LltQpqdPjYN4kFNvGogbEK1XNecR77B0fP3deraX5nSaXy93Geq6o
FbosDB/OqCghOZEzhY1nd0m6BPILhk9xJKzz6hMHxV7aiSwNK8b2bF9aTtoLE87AHG2GtsWOYYQv
eKePyHyN4VCSqoVfXzH7fiOK2AhoavytNKIfzV++z80dnZHqIAu9qtXHhlYFkexKT8vK4bJosen3
6KmG4ZKVUC1GBRgPtqX0S86asYTFQZHknd+FUV8DY7ZVSmvjityNI/6Ny8WLzE1TIQbimR8ZZe5+
FfjD/gu0GQGrCaAVxmwwajKd6RM3BwSIye2X/hGNu0UyObmiigv3OHij2Tj/F77bHCfR3Z3hKuS1
Dr97QcnhMKayIW2SU3Y6JtqA7bqWpu++MH1FYHj2/PSlIuw7N9y3Urir+nEJaAX/CnhtM1w8z3zB
i6LMLRnZxpVpPbunf/qkQwrPG4HpR6mxiMc+VJKEBdX9XM2ugPYSkWcNxRY7mnfabQ8ctBXgYyme
zvs0/tkWV8QYAaYi/YEe0YZXPiBgoUfjmtNO4TD7m0cAGEnHnah91P5LEnkda8QJC2haptYXnrNI
I7AIu0gTZDI5A6AX1Rua3Vc/GHS0U75zQrLx7Oblw40rImOuKPV4OOZsXiAXQK4JkRfedmISeDai
x1sPu/h3Rg92XlovQLFj9Xl9B2B+TspAHh0u8TNtZfS+NVlYYfigCfExpVwuwL0cgVHQFd8RkjRb
V3Yfcvt80XngSuUz5dH048QYI0f6ZwB/MQ8J8XqTKmP6UPei7F/MDJ+130a5ci/S2R06ip8KRyvw
PfuAbXiGeoXqmbtH4JT3/+elEaMp4S/3B0GgDWSnV820HxaS+gW6mqmFI1R1U31g9Qtjokjnvb86
1xNDYF/pOE0pyQlNsL+d7ixA3pixALObfi73h/b3iVj0PBRBInQ33mDQTvGNCltutjTq3HEHXNlc
jc6S9XKYItDWteexLT9Z6fxKaEK6P11tgV0JdB78j9zRDuMpoS049Lwj7kJ8CvDoj1At7LAhzifG
f76616t2DEIUgJJ5EePmHaBLYlb1FgV1a3ksM3GVQ4Y9zwwM47VmiwdwrcHqhv6K6IWNLZAOBSXD
99LMd6oteYsb4Eto+Ewok1EJPSKInSJuVof/l794hGb4FG96JVneRcRXGEbZyvPtMgBED4fCws4D
PQIOcbYfNZXixqCnq0awLWBs6KdNst5k7pL59lgeK96KdANCE1hAf2LL6OrBla5v6+ddNm5f/mf0
FM1gDnpETn2U+gJxW/9Oej/LGKOu/GtcuLvE1NXHYmzIK8NYlpdbKVmFhrTT71lTjDFMKqGhB6U2
Mg4WkIdI0lCN6E8c22XGr2e2sbNWJbPUqxSottwpH2eexOAvVJKnAL6uvlnCQanldj5e1lx+69Ka
9GdOyZTlWPV+eWKbGShx7cYFYgrfkR/P00sVirj64T+0api3QsrfV9nEgipCLRPdhp3mnu/QUDPN
P4C42zi0eM8DwoaXlmxCEebP6AOOy9oNEThx9Yc6ja25pgc3zpzfe80nd5poXQ3jD+q9Pit/YXOp
251sAwrZBALD9kvm707v917C0qLd0pzDdxCMD83uqmnvAg5czkl5iG5+oQa8S0f/2zTxWELrftnH
ExYXnX0dTl8hkotvRpeZGsd9Rn7JZUrBc2SV7Wl1r7uztQPQhbDTgSFz3pnt1v4HPboB/sKEg9bq
YXNUmYJZ4EuIt0kuvaKbhIkeJSrR2RF2bL1rhtfrzL9pHKzZQlk2INK5NJ//PNKsyZHxNeK93SrN
VgXzOpIVMvMBF+7p5UBqQb+qeB8JM6qDvxfHNmvRBD0XV/eLen2TxT7fG/6l4RMKUDLZo/yKwDQJ
cHCzToShRyXhEQgPuc5vzz0crwSmXsFTaWGlfasaBhSU89QDblbI4jDM2QygXmoCm7dLoXw71oDN
YtiyINlQtGzV+NDkBE0A/1/eaF1RvNuddiXOWY/xBI0zRpbWxVVXftVvGvTuMkOIiPkmdydnl8hX
3i/WkifPvD4I7NhainmGzsOjUcTE1kuIzOZQOYoehhO582poPhVzLW0j4vwPOLFrIZYAJ4bguxf8
e4zA0X0GsU7tl5fpCO3mqm1bDNuc0fN/Pg2cR/sbmBJqRORIyBgKdXlZyRNrE1+mFjz1/K5+qzAU
jgVZSgJO4yCvhUrFcaI7TXHBPxNdLgOCdf+aZhW2URhSanDfQSWroHgGBnG4LF1uEMspiOum3afR
iIDl3tzz/ERrUAV5WF5UiRvzKdn/rsXZDh5BomlSFMk4iHgnCI8oNy5W/riOd6Z381tjvInBmAUu
HHHazsGt9WLqgF3fImqfDMsCwladGI1yKlA35VNcSoYJWxzaCQnPPBOiOH6TIJYmbJE2+jAaDPAP
mLQ2TcAicRl4ppCFn8hkYYRJZOoZs4umjrwYatYkSNYyVkxmQAMk+GHbNoDaGJjSNUOrtKkdPRYw
Kbey5Y/vUUEpbQ4F1HFSop5K9PGNIBTvokFKYokkkqw1gfFcUl40cOCxVsiBW8eXDyTikdEFJN8Q
n130L5vpR6TBGlOjpE/l64zLCn3GO7qBplB2u7ZMyRgdfoeTxQ24VCywNGpzQp31/0OxYs8GiwAg
5BThLIQYPRUVoP1bHc3ANSMNyMOTign2NalllwrahoMWIJQR3eQV31yKkkvb4Ly+u2iJZPWbZF6k
UVR2L4FiAn6HnYY8x4fapk8zfFuoG0Yv1xjanDwsKDu1sIHwq6eaLRIt7FydyQuQ27tv210zcEC+
AqmrHa5N87t3Ipv44fiRiSmS9FRtJiX/5SeAPOA0dCHITOSdAZTwWLlwPAditYJ+iPh37uFBg/Jx
mU/4zypSNZVrE1X5zXGgGUoUkSisYjONwlM44Ifeocx+1kDQGSdFx2zdas+5TK42xplIpK4MtKdB
nmDPyq1joDBkb3R2503y/B8a8yqPojpEH372R/o48RUPuhG8SnN0NYkg3PEoiVDoeIvHvkff3I3q
JSlRhO+QKoB04b9vY5Dxvc8rWBfzS4wG/2Wrt9KmXvk6Ex3UcwAxq2z3HqFixLfxvab3fNd1HQhO
X1GJYllM1YK40fmRWzPfDqFxUkZHqNkAlZ7YzezxYBxYjpf46+jj03wImkWwUS9Jn5Z9vFkOvwBJ
K7jisy7o2NfFJvT/rbsrVPxFkIUDRvZyymN+CMDSPI/gYbxJane1OV57zEKhfh7Qnj73v4r4jRZT
ieFrayBJ7ayajOOQSqOk6rdf0t7HMrN60W5UhVFaBRD9KspHANNLiijrBZI/tD8dLgtwRahNfvWx
QjS1DZoitEPE7pXFhbOsPUkI+oh03EbMxfTLgrzYYU9J+R1e6ZJCy51U9eRwkf2gaERt3vLnm96J
+L1DBQJ+V8vkRiKrYAF+wzh+32h2kWT99pMF+NIXzgAyO07mrZq5Ut2YseXOhJtOuGVNLopqC/M8
o0nWqaeQCyWJn2hvgc3DCBB2SP8c2fd9GJSuQj5L1A4okf5hwqXpZ+XK2sYaXeojlbnNx1U/WxSt
ComM8OUjX4gKHjs9QVrhiYRehF+7TgmjSReVssqMOJL13h+mSWEtdNrKccvP0nGKDQsNagIwt2NJ
uY6Xnv+0rtIqudNnRKFne/IqoQKe23emBzfd9Svnhh8LXci34sI1gTyk4HhrhXXfvFqPSQpuQUpU
JGtsvRXjuH5BjZh966ci7QX9/vX+kLVcKkMes81BV2WYhE0zSWHoEv7s+cu/G/4CYxJEjISidI1E
u8fct2vj/UzCzpkirBjoiBrrx9+T2aGP9IkP6p+jPV2/4j1pYexpixt4Ei19z+UBRE6AsjV6PgaA
gqFv7UFzIj3ZS/ur1rlaEIMmJ/t4SVwswkdZva4eb85MpN+ewAmHR/6Nfi+kkmlFSjnGCltT+hkU
jSYuCiRk1q6eoDkvH4js85hUpBKAoFFv+lukIY711SXZiexoOAnNi3px8L2zPN3aDLsYt00EIiAd
GcZ3rC9hXkgPvkPcVMTIRCIkKzybOJ5XoWwkm6SjfzJCC6vtXzVYOlwYiS/Lr9k2SVGqyEFWL9K3
P4PVW3fgaC2ArGQeN8nK1TfoyedcDWZ2GtFDJtZ7IezUxAaUDI4m5xKziX/7gaZAy/cv0lBlFVmM
G5hf+u3z0+xf/krxUeE2GEWVK23hWy4AJNTAh877xWSSX8qlzss4UgMSt9DqlWEdUvhwM1tCCA9m
/nT5QEO9LHe/FpySzH+dOEthL5KIge+fofdeeWPlRVuCKfaTxlKRaqsHcgX47bne2IFMWo/ht5Xn
6dWWy18lPULqC+WrFC1O/U6jmwBgDbA+nHLK9XEepWiVzitvWwf9fSKYxrcn7WsR4ZPVUeriBYa7
KvolCpJZKuf5hQ4FQjja0zoY95v4vtINGqYDG2wQLaK/bSBrfznP9gAalBi7va7FR/kQtI/+7Ssg
QMB39gIIFF5gEUmzPhfwCAXgSsUYbRukiahYvyxtyRQShdPQyfHh0JJJmdvmUV+JChnMiP2aQ2Ks
6Uv502L/xmTEJWw2C7v16rKaYZE1zsSJ0uNo4dYVtjdeqb3m4UvVpfiyTG0lgfWFd7mbuBB1Lg/4
PCIK7ezCpkuL6oo5o8hMM3pL44W4ihLATGuxXMjI57ms0vOdQj9G9d4iCGREDHRQXhR9qXVA+RKa
FqGCFysq3dZxS+yG6ROSls/fpWXzMEIL8XWckuM0E3DHRXikZrIUJHOrKUow23Zx85VW+YvWoVGA
if+xWbT1UF9nbOy6d0HMDmGVuvR91Wm9jSvv21y0WNasmjNKJBxpQHGXy2x9ay1jvJAbHpVXA1f8
lVfhUmtlyi2AOrgiM8H5KsCmW3U8arD6OmaBvDG5i/OSnqMq64aHza9EvAWKDh0XrEd0doBMLj2k
WHJ7qp+WVATSgm9DS/CaMOo2rwZzdRv9Y8zzTpTUXP4b1HrKgY1//kIHOVizcx6Qg6P0HbP/edgY
HkDkAiDijHFmEU0X4aoWR9+o8N02NMZb+GmLArOmFZkwtcgaPPIuZpJe8yFgvRYxUx0gTzJZpVLW
bu/jQrl0lrznQV8/GmuW71CkPbAEsZzweNfdtvAzGdk4phYD284GqC7R8cn9OlSw+EldaHZNSp4n
wh3TQabiBHMjEJrWBznHIlGx+syY8D7vd1A0xA/T7rwpznALEH8Rm+xzTORyRzNdeLfnt3D691hI
W62B3M7wZsS7sO/uWaGvk+pyGgEh0KYZ3cEjsQx8/umjWbLsH5pLSpKTmK0qNc2egngIr7rIqOEY
L6sE3fi+4tkI8cUV8QClzEMAuGPilrCkoPAN9lGXz3isv8prWDnKK1/gcwfpiRcHl9mF7lxSHOEf
M/gswqjo09iDaTW+pU0kGVr5Vv2mItHgr++57f5+E0iW+OICfvSt9ZSgMXdGVSK/eXMNpKUMKV9N
mg0HPrmqk+uYmt6wCX8zP5/R9qiYlL4f9TRKjiMEh6PvePnNweUMCqhDovsp9JyR7kg7NlmZef+u
qvCX6zlTyzMdRvp5lmCvhYc90qBao7InFh6HBvZD/BBtLJzhjgawXc41pR8KkS+HV1PYWjOGVKR9
ytZ65Hl5DHsY4AW3W/rG42wBRu3ZttdlRs8rYpRJuNQTNydkzvegP02BWz3qSwmpvnxC8D3Z5QRx
Y346jSoHeRwMf6L5x+9vbVmbTG4k2VTFt9z+C7KGCvWN/JWLFN9uVr9x5Ak7NXYL189sJdGYsY1w
PWP2UfoyJDIC/7VmbbwygDOFjrM9rQPTrr3ZSUY5/Is+R99IoNp4qNCdY8YetBFQeGoOZAIWxey8
1a8MVNvoVSEHuPqvDmdmcFZD/z0AEt1GEbP3KNARK7vw48hOb47QBn92Fu73fY42Fg1lER2ENM85
PHcsdVXzMqlRqfen3mYUZUQ+ltAsbqAKIV9pFjg14dIKCPeqZKQkFUjXqtDUuNoO8fvYKUJpgWks
vPFORD52k0JANSD+g2Uzpja4lIjW1v9eFlVAzzrb+ny/rsWcdWUOCg1qgxPpOPJ9gd1K7mRJ2jSk
jbUkaWP6OZPWrKxxiFoaUxnW8JZIvlD1JlfCCd+Yr+5QFHag4fBgv5Er5RNAcgmLGjHuttYHSgH2
ytWLJWuSFzeUm05ocFtdJymsdeMrk9CNwubh2LQmdZK1ukYw+euDjuDggs8Y8ykU2oEiz65szKXe
P1IqllGWWrDFj4/YwJlQzN+JS2Ivac8EMJ63iq2iwk71xV70yZ4McBVQJVWplHYIbzVJ++f+ZFPR
5gS7vC3h+oOAc+qGlonTeQU/275rykbQD0AQjDLA88svCcE4BKUB9pOrJWeuAXlo/M8XPg/ACEMd
3TcLkW7hsGT2ZrPXO9mBlK8xbO2wa1+2jF2cUL0bjLJoEW9lDFeq+YSCbt5zp1PPRmDME+QLrPpO
33qKtl59nId34QMMagO+9EOXkUouKSkj7XT+/PSUdtkX4+gwYqaDpBnkgctjVGnino4flAPP9Lu9
HX60nFnF0DPYLp+wLoIjsziOcmusODtaqPfF8WJ+qYib3Kj+MJNHyapNZQRU4MJr+qKFwdYAqWfu
VzjzH9SfPWJndvxTZ2ZHskJjblQlnRjyj01Ql9Z8BqPb5aLEdrave3mf38IgkZDwdfArMi2+tMlN
Gr7ce3XKn3y9Sy3EV2UrNz3fA8BFj0AOV7GzuBZ2O7R/XtDt6Btmr6yfpolrNIkFBjIaOovOB02x
gbV8k/Q2qRR6se5tUbnshC7esTj4f3xWBf+PYiRO2BxDKZshAVaboSSgJl8gvcY2ptK3w/ZCEvtj
/DXWF60zGcK9Smqrlgw+bR4z109dSZ8zLvbdGxaWmjdNzBLHzGqL6lKmltwNLL0wy31tHsyUcwCE
zRAnVVRpExrIUPZ8mMiT9LMWp6qVJVPdxHwwQGS1J/ITQFYyjfRJ1mNZjO8Byn8g4j7GYkbaO8YK
WPXQiHW7PgZg8DxFSjMJsRFvK7OVaAbDvflXvh1JyKDrkzUyAnbz87VLkF+38nEuT/xRTWP6Rx1g
KOQEBx4xLtdn2se7PIxmsSgPoneD2pZZPh2EbxZj32ek+VaLpIgKtRdvtFEz3GdXG3nmsD/vjOIm
flJAQUmGHEU1AxOlLEeUqkEcCGikzM0fIQY1mceWpJoiDdbRp5RmAf89eQmxRFz1HOvXwTaExEzw
kn3+JbDTQLYMrCo/+l5qrx0pua+teWgWf68YzocCLIIpOlPHKPmt3dGCq4GjVj3UWRCKknYYMN8u
ItsbjLuv+/OwDWly6si2RDKxLijc8cHGHhnDXSz9v9dajO5qGKPpIy5YrGjj2OcxqpUzQCOGc6bN
D7e6HSPDOptSM7f279nS4Io68S1ZVZI3uDn38u7CDCU21z7D9+Xz5JzK9lj4rP09dDXZqMuiHFBq
CNMv9hnAjr7QLqdgZghIFgWGRg6m83W9oOGPJyDRxgP+NQ0oXM9TvZwY6unowY5Kp+utGdo8NJKk
usWluIXZqWvzc0TCoLB3w8kQrufhIP4S616AVjkgKnjR3NTW/h/Otitym6+zsc9vUqsERK3ebMMr
eyOQJnHNlMwFEJPtUtaujYwSrCqBqgIkkSliEpXFESyj6pV3gF0TAMWBJ6j1lKapbyApoyYBVrhS
jOdRYHm9rExrl/G4C/EKFTkokXRmK6bCM/14g6etHwMjtTpOP1COvH5oAXDjwwa+gpRa3k1USrqG
YLLswETW5BBzd7Xh52u/n2w2XlHPqmJ1uz7TZJXBRq1bH5bFYzbRKL8OZv/zPkNfg0ex1buSUTkE
Tvt12UYDxGX8Ymg+BwRy3VLgoGq6oaEETnZPRrjUIDR4LCakAaebxhGtcbYeiZwz5dNlr6hQgQzU
0XEnWnIG4Cj02MLjZLoYdNX/UYQC+D8gDr6hh+mYer/q7tbMIcbYZDi+82GDnTgNdRxoJrVs42Jb
4OyNTiKOZyj18n8wyxoJLN+446cu9+PVmaFhUAibGCHoQVDV9wXxo6+4yV+rafpnugwwtTqPIqGP
hHOOpL9Wdq/OVcyxLEUcyktmcr1ytn533qVcWcTpZYvIAmjq6oQze9zqqlmW8rDJei2KrCk0cSz6
y2pbX1KrDa/NUiUrpkyUhlL3ZvbpYF3nXG7HpNIcYoAN6YFGW8SLMARCgdpeJvYFrW0Sj8iuL0Bj
iiqu5WbVH8WeohTIfq5qAb7sFstOcvktaELUiKe2z/IOfrK8Gm88PaRrt+PLM4rCn1REb0ubEN18
qv+Wqtx+nE4BqoR8PWkty1r2iRK3sSGLquUTaPhsXF16LEv2v0nxAL+cwJnjtuTOPFLC/t1fVoaW
E6d0VhgYtm1KzPMd5J4NXMginb4mygcvXzaAdT+YqY3c4vnn0buMxonFWdu/ho8FvLVnHitJjlD1
zaV1NN54AtlniKi0NDy6jutwLNCMYOLs1YxTxnYwcbrzhc7nhWBL28Pqa48OR76WSFfDLA4DENYr
MYTzEejqsY6sXSuvY3ezTkcNQ2zkR1YOT5pSM7N6BDF9CK4sFst0sUTVFGxhL4KJV69A0kbep9vN
5dQ3sTMwDvp4iXFS5TJTPHZ2EdVcZ8mmxTrR9rI2+cKHu7WnmaUOTMAB3pz8TsAPpR7TTn6bFOZQ
qfpCaMsu236F5WBwO3PjBVJHNcVTehGlcyvCeyCg033tGggvgzVJt9Gpzoc1GsWlqrkOLPn6Lc7k
GCii6uxCDcDTA4wMbXqCb+y4IZjBRnOl5/PKoDXka6KtWwQeMzFZuAsWE0RSd1g7h2xBPqkhpgM+
pf/Flg7lZGeeuVl5Otzb5wGYCF58B6+I8V1jYBfoin9J9XBI0i1jBmxBHh9AffZ2hl57hNCIa4BW
1R441ltB1S3pMHCEi7HJMU9Ee0s5V+YmD7+QhVa3HWNSgm8lOAbo9JmhCPcGP8XeLnKvZWJ8Rvvk
PL/l7zVXix497EjvyrHDbgo7muCctPaSBoTNhokjMO1qpCrwRwBym7eDicBGLD7yzC/ND/tT2LfZ
xCKa7HKltIckgc0nnS0XXwWwndw92qX0iCzFuXUR4LbJb8anGnCoCgkOamMiS/oaEA+uQAKUW2R1
BSfy1cFihsnMcSFSG5ANNVyIkALK3M1BDk5PqaFohHLREAGphu4LbFSCcViWj2ReeYcZi2Nktfpe
v6s8N/yT2yAAqWivLu+iNbQyjtbN3KThytYSjySG2zCAzc3NHdGkt6X0xqncfpLByFmyfNHFFUkK
pu1JIUN3QCyfRBXnyqygglOhzl044pyEI+2WXoBvOdhrK+eEOu147PF9J0L26RDL3yyOEXwjKU4w
8t28Ytl132Lzy446VyEG7YJDyvXtnApG5FStmP/zznrsj8vWq3F75jJOfZjHLXUox269Am9g1eVc
uU0MNlku3s09+HO5ihbKM8sdz5FvPswWJHkcM9yYeaID4MXa0vxc/qslfBf1rBD5g5XN/YXo2gKi
aV/XF4lMBAcJiDxwJG7up6O0sdKwoH47w5uh4872TVKsfCBaForovxtmWMu1rWoCvsQzkYSOk+5L
kKr+9EmeBDbwd3Pb5HX85OGmr+86o+HxtIIGnRkPqif9rBTvpCMNPzs4L8iX1ZPt06Og8fTO+Ilc
Tafz6ZYMjmNzdvdEe6g/ppFLP0IPul5xIu9axkIuLHXwHjdZwH7JhvmUjbR8iUpXP8n3G2YtZvDV
W1qR+32sg7mhWihhTcLroCxNngSsQ644hciO58akLFeb/GbbA6JcAOAA2596WKJmPmCODv/12MzN
h378HvfJkfruiK3ddoaNuFb+uEexBQDRbbvq3z1DU3jqoZF4thDCTSyst/wn3RQZRkItm+N9U4fs
ahUhTScfEL1oKNYjOZPe81UHzUjzdE2QqSo8OEcGz27Q/ayP/BrGqdas0MA6Qs9M9cUGnQIBPeYh
HSFQqtwRjDyabrPTWkdCpL/xE3Xdu2elISq6penyuLGVPeeWzZpPGloeXIW2h87fVVWv8i9hA1qO
slU/hx6JqNm44OWtOayTvurHa5ZSpqzMvXRP+bdO97qTuw215vUeFHh8OMa9rUyqHOiNq5Y0CP9z
yvnc46JjSbMjjfGKpETV0o27qfvyOtuM34rZSLsDXPiYio2d5vJrw//rjcTaky6bMl1SDD1tg24J
Js7D9rr7Xo3F2Yvb6R6o+Xx9pWaFzWqfDHv4kmjunF+EB011y+GQzElCIfZNrKRgwaulD3owo8Ot
le88ou8RyplZIADoZxorQmxU3WnrdSZhxxwYFLfnz45GhLr18vClxCyVReV+3WEaMlz0njIuS7PF
Rnzm7qKo4s+0fl+nI8PfXYbdqujTCqwGgoG4hAq9w5H01Bj5TsCVSL1OW4SnC7Cm4Hm4BHRdroz0
82Mn5SZ22Twb4F+/bkUiJDH2NYfoxyTR1ulRzpDVFtk3E3FRrhdWVdFPipJfC40izyhoFsDljhvO
aOElSmIsAs1rmIZWfBBN49hClZ5O+9NF+e0tYM+8HWNHeVkuvGf0MppX/k5bpz7rAnOYGW1wDVRt
wNrxxoK4+xak/Stkp6DeJbom5DXsxNh6ZcPZlESWmu5d0T5tfkhuhzLsDN0VIE7Udr/V1zicnQLA
MyHnnEKQnzRNctunNIyrcSF5auEeh61zacR/bLdTwgiayZcJ3LofCZCWjmWhPSZMFwisZqCYJxdt
cF2lpXBMPGN5G8M49mjYX4xDVkBbyMRsAFx11o04h9GbZuyUkdHdkgrwFOyOHAtpdGZ5cRY7sM2U
MmEhfOUC1E9TeRnrfVfLhe7uZpC8toesC+pY+vBW3bAtVu1hS05j/i0M9PJL/rR23dUQqaifWatq
s2yYF4IEa3wks1gLPvR9fnARsztYfuWZekEQqoZXcZ9ntNspa2SMaHKEEwYBQQ5Z6hJAVg6AnNbn
AhlSDxsrtnhJfCzMrbxGqfaTf9OzXEtLGGeMazGMGWSVFxCfFDQoZLg7LDp6jMY7QDhQftZT2oYJ
TG+3c3CuV0h55dEpKr0jceTgvxdWbzWKk4FwnfEpsqglOxGs3TbWiBJ0z3Sxl/wimwUYCuZVcns+
pFIR/9wmq5c7F2Vde1CWysZgYaDSYIa2gd7vstIfCnkJ+VtU/7+rZ2TcySl7S44HnXWcGLOGLlcp
aODVN4nq7D+7V17FEhcz/cJ9V0njD4YXS01q7VVvD+MIYsWm7lccuwUgcrfHe3QczTatTHjmVFaX
4u9SFCjuwcZzE/xxKGRRFCETVrcbpXot2aOhMWRQ3jp4KsrWcssNxlYdMvFfH4aUpMM/cPnupXS8
BeI4yqVlAJCrWG23YHPyOfKYMwVKz1cIc7ZLqEW8aB/aKUrVjqhCHc/A/H9xwlxUJvwc90GGQU0X
DVPbK2TsT56bw5EIPElWF+3Je3OcUNlorXPLW79ltJ2b04m8RIPhNRkpr1L9SuTT5bXqx90Wb7JZ
0gRvjP62z7MtGisqJx3WkWlMmEb3hskvsXVBkq3TNDeCcgT6wsq5PlywnB9qbVlS8ryrIj2YFZ+l
8b6E1TFqkTXtG3pkdq11tVpSFcu/5UYuYIHdvEhVco/pt0XftkvDaeYR3fyEZzBXfmJsFVVDgede
yD3U4CnoC5NOzo+N5Py0JilRt6vMO9pjUkWmEOlS9CZ6CNqdGlGZoFQZmt+eJygAFsZzGm9zTC84
oPcfnoazh51pCqFE6cgy4nFlZbMcZZlCW0ANnD98Cp6tl+i/mqZ+ptqXII2kZlrrJWrOYgWlM+Sr
zkxy45QgOKBqx0SMPXkjaYB9KeHzepfEzbDo6h9kcCBJSC2rnf/izLl8WayNBy7a+wyqN1vD4tmq
pqrg7IoGJNvXEOCJlkjRH18nPQq2MG/6Vp/sbjmB5xWIuOi9ncQnPsbP9Md3dlnOS+64ppCk4jmt
Z87A7K4hRoUxsFJUTjN6eZUoONb44o0h55dbIySLqNUZiUGfNwyxcq/4O2dKMw2i3XDzijvjtCVm
bSQxowYW7jgeszkmHh//2KzAbUfTBMF1zuGP2j6K5hPOE1LO6IQVaIo+5xjuQnbiH6DLpVeup5a6
V6AFW4w+I17i83iEZ0p9D6adfetPCTj0OwwUY2loHtxbFKiWQTl8E9GFK4WBc6DlZLwy/m4xHkwE
zxA9jlSEFwS+RxxZl7cxDdNUZc/X5lI0nxATlmJBFPKLKxm9w4WyEWM89AdkfviMgdIGJ1BW2bV6
tVMIQn6/pwn8s74Rl0oMUtOwamqqmuUrlUyA6LP/1nSlROtNIB2AOctp1/cNMf6bF1rzUAWj5YHG
225KRt0YSkwWuNk4nqm4fAoJC57GcKFAhYhuLFCFOXGQjOWJJ+M/W1RLUSmTEqvJjnldiOxnU7PJ
mlADHHkBYXw+j7vrQhNJP07y3hni6XJ+SaECxOD5KiS2ab08U00ILU42QFweMWgUrnX7+IL4QXRx
Md4kr604Ru3v+4PlREDYRLnt+6RHVBczD4Cb8RjX4eGxqHF53WUFl18GNdJ0XCKkT//qwfHbC31L
XgJhd1sGUkl8+w25U84rgwjgvPUBiAzTubPXJwnUs7kWzK1Yb9ckhZvjqeRjmwSYGYDHkNO5kFpG
44WwglFWna6KcNerCqBd+HNnKXDjxJk7FZ3FWVda+cKhrUuiH4mE8dAozTRsRRVzl+pPC4EBW3Vs
WAzE2t7eje9jfjh77Y0w4iqqIMZQ1wvOQNq6EewxsQ7pAOvUcaw5QnU/x+pXxnw/2qNY+Ek7+tY4
FZoT2BC9MgK1T5WQWX37CRQODJu7bpQYflgaAaW49gKE2WxJIoxhyjkbcYG1stTmsiHjULPctlCw
j2rKU3dgwc4S6h3CFhojLXG6kLmz+KFRGqxPqUDzlGjqzsOqpFCPZwKsLV7Ak5D95Jm+bi1dMkdR
kSml3Ne0LHemnrXpn04HJbRvbOVZWZCCOTz4mEVeydzD9PLw3MMoav6xm1/O8a4Z5wSZZZ37rlHj
7A1WwHTpH4otqbu48hIUw4K/EyRYuwZ+ZIXHROjisobwZs4V68vQc+pQqbhz8jE6fB+WWgARTLMV
KB9FYLsPiFeQerz4+e2VT/ZPY0nDurP4QPytEumkaBf9RJJavUVuzcQvq9fL5ruElVCZgWzxc4Gd
uUWH5AkQIzk1wI9eRSfeiNXnSwhOm8gCI3tyN7Us/UsoHQZiVD6Z9kmPIvUhm0Yg0lcbRSeqfvVD
uzm7AKCnw4KhASmTlFbYIZmTFljZUdb1HDfbZoElBLGCTReXz7aCkfAscj2C+7ts+gvqZS9UK0Nb
29FXc5us0TsNJM3UZ6NrsgNlLCoYQVwSm5Yyxq0STmJWDdHKhJ4pK1VyRFTsenGRdTLBZMqM0GB5
WPOACy7PzaBs8Veqrc0u8GkX2K0hwGPflA74W07B7y1Lkkf3lOCs8PTYPmEIvAhowMcv/oZHKl3i
rXq6/sGJh+BBlH48RYUsXM2v0j6fB94tuchI6GZDPNEmoR66ECd9Z0BMqA1G+Y6B7Bjl6Qy/VYXN
716RHoeNaxAXOXZA+QkrsnotCEnA1fdQPHWPZFueLDBbFmN4jiWAuPVMto2W03xjpq4PycnZjXhB
vqWYJ2taZUTrvvzjdiIFhf/I9OAFIo5qW35TmwdoE6MxjvcoIZ8UUoaUlBfv9oWIFylyA+Rm9Z3H
XCglsynulzRvZXQ29IXO9d/xSNcf3fqZtVP4Bq0mZ0MycgE/hCcsQtmaOKyr9pQqKH9ZYoePRg03
zaSnCzwEV5yFyMj/ir4UVfKXazrqgi+k5xaz3tbHYGcrfGKOVAx8R47sxmkK3PvMSQ4uSCnsgkAS
aRkfTmNkpugpHF3tr8zvIanjmWaa5uaKCN9OGiQRhjlzIyVJv0MMYK78n95wSIdp8PHSHHYkj/2t
vVV/wOZV4HXaoGmEeRnwvgZ3djzKFpqvkH41OdzvShm3kDpDeQXID2NVmUAwU4wcgK53zdHoTLEW
ytl4K61KFzFBqHtGiHMKkn/nIDhiKlXC17lpvHscfsQYaxPhYqeh2aE48hOuaDrJXAE2deIAVl72
qrd/h0UOK450dGST92nSnb/coTmwZ5zjiXi/ibgboXSJPsWWAjthBrpXaNR6OkCDmBTjAo295iTd
kSzaJAvk/Tu35PMgxJ3PNqsZiuYVO4glix9aqbg4SFUwzHbdP7l9j9YKqy/THLjxPTNu0egmQ23f
rp/pZqlA3aeOPj+E3ERPb/Rfv+2ADcEsq8ALjUk7RR4zZ4MAhFUMJO5JWykDVBpZONA8o7r3ynWr
ayzNBSalONYLOaJf3PfdWRd+PGjXjkXefV3GEEkNtlutOLPNfOAO3nOxbDX87+wdd6xQL/QKKFh/
eJVRlJD/fpwFAclGSPgazyQ7YYqBnRBfdP3G6kLa3EQU14f6uUfXnUk4z2llQdcY8HePEecYow8f
sCe2X4kQN7KxZZpZeOggf9UOc2r6rkVtHEj+wSqs20Qgayaezad2QcVRWW362lyXG7SPF8JVUrDI
jGZs9JYNAX6qnTu08OTow1hFaKY+tRwz02pg1T+sbf7UYHHMjUKykiWfRbwvkIR0NH7fNTXU/DdL
PGT5eBD7qDBJ3OS5SLRrtw4S8YRp0F1lhpXNHx8gQh2EK3k/fOMTr+cuUjAvzQ46Nkjg/9Dxwa16
WozenYQoRel77fGifOj1h567El7L3FAktvyRS2BKDi+9MtnC60WOmz9mKj0BS+mG6+V7vUmKh9Cv
XU4nr8IsopWuNlnCrhNA0IdYxPcUsYUI7jAEcg3wE3RKll3EehkaFFb+PtFkOHAEU4fB9m19L4Nq
qcuxDuIu8s+UxLhryTVrUGOvzv600C7tH1IeKUEaAraKukAjscHpVS66MKNPb8p51UyI/Y8h37Jn
Xb94NeEzGn5CDSCuwOeed/oIM84aF1V1uu/39aozySwau43PoQ4TxmfF+vLaG8ZYlSt20E/qZJRb
buH+IadDGi26B4eqJFWxgdz4xePvbPvwkDpaIW0xlcF1uxpQp5pXgLCjrE9mG8qmCaUzICCvFfCm
OIbbnbpqLz6N/05FlnIPvYsxFyLxzSBA5qt6nS99+B3zT7neDHYZU2/37+y547+EQ0GIHlq9PWP0
CL1wtnjgEMmCKQsWxx2g7IeSBNbBd3t9SRxb1RRFtx7avRn3vQ9+bQr5kGQP+QKwSM9wUDvsskR6
vQV1RZH2VE+HyQ+l6nbR+lyRx1JcyDcNOaVFxQFFrrIlBEH5TRFTtduI6gQ8A12s6z4VYp6B2gq8
+3xkDp8g4V075daSZOn7AJYMZLluqvBh9uzLTqsR16qZN33x7Wpj22Kpg3Kh9wTB+Z7FS75FA0T0
qIfRbxonsFuVm5wXrbD6xyLKr1pODlXZBc7fSNWrOPtE7AbQdWNMtqQEIUw7/4jBnXgnihPGKMkZ
gxn+xPsrRKIiziY5Zfej9GFcicEXEBPBkf16PUOpQ4ktGeKXRm0TrPPY/F3n/KBGm4tiN/jCXozs
OsfjbwrIwB8Ys+8jqr5jF2RSmiRWvX8yhbV7RBp/mZXXqRAlEK7awrREdNU6w52d74m0IYF0cJSD
MuZpxATjmI631HxUcr8DPHdxVHF0X1d7g0mhupfpgvNtYnBay4xuQ77BSB5MVYuu4CbJAyhEhYAS
M93Vab4D4HQCZayevJHdyJ2wpHC9/9Dvo3zlQDoX62UMrg7kbNpFSirwc7jJdzP6OY0EMOqaOQ9c
qGumqZBaKSQMr4V6pAsTUfvZ+ovis/BgDOaaEuLGqM3wDOvcpnQgj1JX10netD6POUskfAbVWDdC
mLfId69AQjF2opZtgrF+rZqPo3N+HoDvZZzAaGrY1zxxwUoBmoXVoQHKc8c+k+CMwijSpThx1XEF
cbVgOfx142MEXMqT/CWFYwMro69iIMstdLnIbVDDmaBRiD3iNuCdw+IzulsY2xbn5ZS+ZsXQ3ojv
+uZglX36CLzmCKdETHYmVuaxquKKXj6f4Uk32OXBtnD9pqTvJ378L7fjBEIjtNNpMi3odGkG1rbT
Z74TZGeUln+rUOphx68BKF/s6VlHWuzjpHXJZ/1hFfrG2QlkogKhwggT1iPYT/G88z+kVrk+0xUr
23WkVlC/evxohqvHZtnz4qLDQP+3TZR6eVwmfc4CUg8P6kqm231doX9M5u6NTMQKQkJ3N/nJPBVb
bYu7JCIrJgBkfPG6uBnd6AmHuxi74yCSTW7Pk+uT0qoyaYs+9sqUwEa8AtegAe0zAToWx7f6ofxj
NSS0ibtcj3+38Mky3kc6y9YKtpokz0+7QOq+qfvrMVRVIfnzIfvLFvYcm8JGe49+pxrrTRG6uyaR
+Em7Xig2rWWbPoKFjihDfBHcbbt329tp0Td0pzTKxTiCncPAf7fQk3+EHR7dN/O1UIJ06uG+QxF9
15olBKvnMkhXdegcY4uCsVFa5hJjIxHlBQg30pKkjxsBV08DADba+04BOfUvJwo3rn/DTlHFKjBj
IvUwjUcSYx7Gak3w7SZOBYCXLWD7jNfzx54tt+5fUVwgVcCYLXUaIbjba6giavTk6RzRllBzme1x
BN/06lnHdod7V7oNp9XkK5tM5UmlHe6ySqP2EajsAjPcoPkjL8a2aoWUruC3g/8ShF+kVvRPs1V+
w8E/BAMzQwK/awX0yOA3ZtbjTJEb8UehnCA7rgEaxak55xdeNzq7EpVjAhDs68XhmFQQ5FGmEfDl
92xx8+xXhLBvpqy7s6qdTTY0JYJ9l9KMvUXsmXEPhcQVhmLapc41XfRxAkseAp6yJCsK/oXH4Ren
tiEx5m4V1gkaI2kivNfGUi+3xwgY7Yyy/SA5ow93SJ0/oQ/qQJ4drQ7HVe6iRp61lZmPVkB4xSfD
5ZLmQuDi4gnmAXc/LjHb1qZouCmL5YrUNQGaSX2SCpBazBmtrc+CKyWLZdzHOKLusR+Cst+doluh
D7F9//uKDIsikfvD0RCSLoXxyDetgRYPuXSsTNbltlNRbzAp71NHibdNHkOHQWbtPs/vvd9ZrVwj
e/Uif+Z69dFEspsxa6A1rclkR3EeW7YyEyZpftKUb7513pcR6qpLJiT9L5RXy3aIA+Wmw5QlBv+v
rBAz45G5+zd7tomNB9naG7nQRamS3j8DKVMLOSwTBztQIca7iSKIeFmdHLDBn3uAknucNi6hkWa8
GHpAlr3mJ8miBjGDSF6YtAZm1WFrTUkbLJlITqOTFoJD12Tg1SJStsjQNGSrZGef9Y/n5oXpXQAd
hzrndtbGoQT148W1qn/+Z3XtgWuTlybEdItoZO6VCFnVpRExipevZ8zdmZOBalkmCS5RdywnRqB+
+rb+ZWI5UjKRF32nB5OXhTjQ6PCnYTEmPbr/9yZVYiKv4Z+pUA72NcmWYDT1m+E+LDkr1vM7q4RW
30eNg8PxQZDv4yNctF35f2zT113hC9fwEpmVxI7DIKB5mqrB2trbaZ69xqi01XCz9m/Ct6UKIBox
Fw80IDg1i4ar79IxOXFj6P9v0mdR8gO8sDKg4Ympi7X80eCHZkkgv+kQj/I7K/Nz1r67PJqJoZWs
JaLEB0BjmLDoDttNzEitkQbQnN4RgzQ7fEnhLqZL8/XCZKGFm3/KdECzst7oqZ8Dtz1FERWJCWuB
uJUTUaMT5ulLBCoK40UM8JxLnakxHEcr2V7IiNd4X+7aW9CHS6iczZeoJH/S3baFg7a8T1fOzIvL
Arre3GitnznLTytkpBKkhovacMlSad1RsXoExAUM9ywGJgG8vk7yDGzKoydhpFFEFiQrRjnSfR4R
zDczzMEViX/gV9mrHlTogpNV6C8ZJpdtDeEyxhrPbQWufQsQa83FVOiFP2aV5ornmEnYdqMFRqHT
oEf05sz9ToF414pDK3iwkc7EltFj7hXYbbpswC3K572D3vwJftSKMRvs2BbmlOqMP94kjD5MuWQm
4/Mdwe2keSTzRw5p7YlikyTxDy18R59TbQVa5Ll7Mc6ECWSdD68O9fV3qepqd6ZV8FG1Vot+EIhA
PLghWTr1ZioROGDpsqEdgI33NYuW3Qo7TZJ3KyJYykmgF5xoHHaNMZIZzLUvmWU63QZHmxd0IqEr
cCpH0yjKekb6B28paZWZi0RFhqkTYisJaBdUnLQirPj3oxDOJ966cYc8lUJr0cEc/qG6iGaJqT3/
PMp7qyMRA500falIxl12jgBUG5ytco3j8nbWCixhHXBCX3srtwQ1L4PlO6lXj9AE6VfDxOTAZnma
1L0Bgz8/47yRy4F+OvoJjStsW3dUL9zpsuaD8V0WySKdeiaDbca0fVlKyUIDRVIXNbunnWnzvP2K
aikcxPsbGrotHM9xWrF70IZASMXvIG1aMq/I+/k7hSJRj+t8Wx546W5+1vJXOZ7jW/Ztzzz1Fi1N
HPTc3OSRXvhwY/j6RE4nHGbJ7A6IKnvXuavKL0319DqDNnNmKjzC/UgxQrdlgBzih8/gdgnBgKcJ
fWa6CefxGt4yjyCrOHdL4ynZ41hSBUfuweQoWUZqmJhKqWjEDV86uXjnWPnsGTg+uFufB1TdNwg6
6CupdWXPywZusOg28k8YQWm3s1EaR/DLPqYuMpDD9rJR1l0Tdb8wXUK3ndnbAYGedg3H30XEOiCB
kqGZO58RNfuPXS8TfzcDWP5dS8V32DGrAugVPhWeWadikyijOzZCmzKLb2KZielXS0QAmwyYpqV4
LIQeh4ZuPsEaDtG6HLvT+WyM/Ipl1RtO7SA7JIK44+AB1XNwCDlG63UJcYFn8PFs6abvHp6X8Okg
xYuX2lKYbPstj5u5QTdpAeIwMayg5Gtf6JTgUMNylXhH6ibi/DRHZwChSxODWx/mMXOEegNIi+uN
mDJ84bSOPwfipipcZoNRmNNAeIufCVDiiHb39NBuCVoXBGope8wxCXqZY2B4MUq+zDdNHkQrDrwc
dpSlnhAs2LJgjH4ovMMmcEy++jO4yzNwBLUlGPpQFcC3Axyb461QsMiCYlHF60QIcp/FpycMVf8t
V2FfYDfDQpRwpf4Fsed9Zs4TqsfLOog5IUmPLvSNPK1SEky+yhN1WPo28XXI/cn5GU7W1PDX3CEk
w5L/P9dVpr8j/W9/9NeZ06/HQYW7LPA9IFByDPkvukiQ1aYsKac6YRZWPGHoDpEsZlOfxTivedc2
c72ZDKIPKspAIOjMdCkJUdQTZGqlbzVvwPkX1gFCK/chLSaosaJByWSnQqfUQ1nJ/xkkngDLricL
5aBT91RPxeRpS519cZ0acqEH4r1QBeETfPB0y0Dh2BFzlqvKXTHP016y11GBJL+aZqtUKOo9k5AY
N1tzZu1gNaxN5dj82CbLFoX5G63zGkYxira61Hz8hUgFpDNzqDOd2Kv1lxlzq2IP5jT9rxrSAky/
rT3633zfxRL0XDPiskGbIROIZdk6RVknJVoWZbi9/9pmhIpNwIGchI785lAFjZNP0wYSHrN1vOxg
8HL7kiBKN8tD5W53xkFY/DSxk5WAXlg81E9YSdaSA2wmzllTn/CSzqx5UQOncgP++lUk+hc4+5uJ
quDbP0MhMtFxX+os0KWUxR+SCSwfzJJaiMQ9GiS1uPhVeDgZMPAZ2se278Y6fqhPwV0O2Ec6B/M6
9kPIjhBJ/L6MFYwD+1ZvVyR240PZBuEDydKUNAU3EbV6Sy6f63X9Uzv66CrqZ9E7US2OZo00yZFC
SyyWXQpzUAxRW/OakMVq625olh0mYvfbOqHF4pL4wC6WEXtmTSU6ImO73pOBeEZzy8aE67f5wcFU
VeVHIW6+4X/isor0LwLYzVtut77becR7zQrimyafsPnOqNg+lIza65QuXey2smiNwLYkC522lsnm
e1XllvokpwE2bHSsDPx6eh2dAfaL5ZDJqO/dtD9kcVNAAALWEoYr4hFJKMGUXxSchaJ1nBs/zIxT
BjEWRcPr26xqPciS27+15P5ndVw/wrZaANOhUl2qBK9QrPPzZGaASOjvLVvgOVggMQrawu7bCYxO
EUHMR3urvE25QNW24L9WJ0yQ1zXvXwK5Ovw544KoupTIBJFgdm1tt0c6yHUxbp6AJJi1SEXogGCi
b57wWPtqMEd1Z4sT9ssTT0e9SIDDrt0CkUgTodaFlbVe33uqWD0qQFGct8KeyCS/AxEdmV+AwSgu
azqLzUcQ+VLE0oKfAqpuWJmibVoRKzwRUZcMq0A0/WjQdMQPjUXg6CBglwNz1G5Lg3kkUBVxzs0Q
NwtzjwKkd3jMIgI45/sXQlokR0zr4BiLQw0JpYucV56gv9eKCAMXZKvy14mvgpUslO2acZrUSEul
gaOYrH12WB57Ue0Ov3eyVU4cxSi24PTsqr7Wqqm7lZwZXBBcdLq+8dRvyDMd61YwjfVsZ/bltQLI
tXFqTEuxl3QB3DBOn2aZ6IvVDmyqywahROUpW9YfkuY+dj8wLHQ6wicg2Pdm28VbQ+A/J0L6mZra
sAcrjfbFxWrcoqtYV/cLuzTa90xWZabdmza1awALi2Tcf/biE0ia/pmnBXrOHoYry9FODg8+7oDt
ptKooCViaRjDWuqgDaakzHowzb81aiufNDhXby+9SlirwcnvolO2WhE2X1TO94EW2p148f4vJaF6
kYB0EV2ezhZ3LxiH0FiQfoAXke5hfrERHL1w2m0NEzYOtfi80sbpcFEq3EWG80DH13b7I2LU8bUq
CQg4us5l4C4nH8Ww5+E2Tw5EizGqoyKB7nVzB46hr0gmjfH7emujOqdPA9aeq0eNTbw8PYU9UMY9
zgiUlghht8iILArxM2KPb0fBVBsw5pYgnsdNakYGdtAfvmtzmuryhxMtHWTAa9EgnnfysfwB41pn
WnsK0TIY7EeUOzvnHYP9IkCdOWexVshSkVIdQjOsL1kpFxEHbPwxebfxBwObSnaMcPJmxfkc4ydA
rAZXK8DoF1GThuiNSBSeATvN9HZYJV1ArGcP0820J09j2WrY0OWw55cHUnNycQhTMbzi7CHqdReI
gJoCgwTzhE95B0JYmqboC3jpw7+ykz3WTkllxy8jVVTyaEK1q4MQsU9vADYtAgHG2Wi7gQbCxq7S
jAbnFYC+bovoXNZgU0X9ULr9UYUCbCir31AeKWDQrXrJHdzI0KrcAcN/8P0LpJAEV9DfDXxaJl81
7gZncvKI31EYXN6TbgLUu9gzz7hwQ2z9AiKBrW8Az/GltO9Wb82L1YMRqfU2VD+mQhRRBfcQ9lIs
qF7cHJYayJyimm66acmT559emGITr6Tldf9pPBsP+gD68RM+4y6izD5+bBpgmuMYejP9LzBOQqQB
09wA4wIKME5eLHacAkONqeBn8b5vxGaTjDFxvl1sLK3C61x+cz5ktJQZ/0lgGr23I1iNQ2a/gsGe
AWkmTJpRAD1iW3qvsFIhW0pQ8WyDy2PjcShsbkcjOuyXgiPaoJuIAIOYpEh1O0rU9sqCRWFcxyHB
8CZUekJENF8qVO31F3GxiDkq5Du+/iaWHrwueLPxoKkoxIf/iMlZX+6fOgIVsnfLnZug59YQrnPm
nDULyfA8rFcsM2IVXDsV+pbOkSlBbTDSeo47E+VCrs4Wti2W0h8BRlqzKgSa1C7mv5n2bFeZs9os
SniXMVhjggWdOQArXxdWwGF61E1fBkEM4dyGVe3Z57A0X6ggT2PByAFEaxSJ3BiITpfV+DT5Irha
5gpsPm0tEn/S4iIdAP+NYKYxag7P7rbME6I8FOJxKD8xaXJBOjPx7Fvp+Fku4frOfGfAlmiXinSU
dwj+VoDC9W/+PCI4ZjrITalts5h3ofSNsPsov4VjXGxFt9FM6Lf/Rs1hJ9PT3sP43La1huGl6OmO
OKGVHRHNDkBaP50Yuc94M5cM3CpIDc8hW768tag4a2tB9IREeqF7D3S6ipg1LiraOeUBmNEtD6LV
scSJpJ5NaDDOilrsuZaiXRNEHid12riR/t6a+AHEwyXj9cg6faL+BEOIh8gPHeFhPxtRqa3SEGp0
9pnrkSgWOT8yCRf0AiEabWf6xIrdJujYUMybmGMQsK4m9Pe9UZvTnVKGzFeGjjxPclClJ7veeorU
G6ljy/LDBBp/NaVWvQKpyMEgd1FeIX8WH6reAPytSYQ6wca6HqF5KNo20M1MT+CCD6EZHHOeRC9f
v2ygHyLk0zQPkfB0jr6IXciVnaH+ST4BHQIkx37gJN3kXyZbeyk/G/BM/1JUKKw4CS8gb1OK7SFP
MZ8FHX1lHOmxS3X8AamEMFv8bnIRLrPHK/CSVCwbJU1rD33cTOip0/nwJzJ0cs6+H7sKAvaecewg
JMADEEiAF3EByvDwOeII9dfcRJp3wTDmiVS6wXNnzqzVWZfKc5QMpdscECruWJiEIbOeyJj+KFua
s3ZZdvYzmnGEALDNsRn4mOUopOdVWTy8cMTurPC4AAAwdnHyWUSN+xw6ywTX66/RATe8RQvX7HMW
i7axFlFqM2C5JYUiEtT5Tkl99x33weEsalbfJMAY7zw/qtk9V3n4K/+vukFHZC1hLf3G1m6FkHym
TiVF+0Do+uC7+ixP2UEYeP/qY8mZLPHEb6ip0XselgG4eDnz/csbHT6kZTdWAJSIbpMVHdWos5jc
VxYK+vORuy3PszJUJG+SjDsUSnjYToLvhgeftce8kg74lUotDnp4/4vMUkwjQvaUpTRwf3EQfory
VNjpW2RsWvc+PaLFOfLeOKVT1S8npynytHBwDdFhhRmt2EhZ5JtOuk3hLfWwYV36X0nmyE0xJ960
GcWICJHiEyhPbzSXJOR/oFUB/2iz3VBaoVLkaOrbZ3jJjs+G6yhqeA9DnCVmIZeX1f3AZgShJ9fS
vp8yy5eTQoDeKbFAvG3pSAs1EkjpOrKQGqqGL+zy2OrTUhWxJY7eknGdhFhMBa4PpXAqvIM5ejhb
QLEp37pc5XSIDk3YZauFUEVPoFQRWTthluSL4yJwFlccMXAeceRpzJBRE5ybtPGy3LBrydMuR4+0
8sQnwXSf20L75wAo6TO3EPSJV2QPwkdwHhocuHkxdnNodoX/KtDJz6cH8hKWqOoUtxPilfv1kO3m
UIAZEFDgcB68DYkJQLjYArPWuOtjlZMU/B/DwJPVCqL75b1246LtJa1albA0UogaIZux/GEwKTLw
6kDYgBjXMl+aI06b8GNcmU/5+X05rqWBVQCjelg7b94Zwm0FrCRY//glolCPgCRKvI8X0kQVFHFW
pTtQCp+fX6bKXy0Cpuj2u+ErROkjPK2gUCfRyusvjERJgEEK3QQQzb9lYPBypyWQotsz5r5sLTz2
ePU5fHoSeKTuCfPTF6r5nkvXkaJohYIwNgiRn9Ma2tw8Z0v4dRuMSOsMthUmhbY5Z9UNLUO5baxU
DvieaWPe6hF37zqewypluuYUwJdST2rMyR/M3ZIba9JAh2CZBJtkygH8+mo8Vs/4H0C9A9q30glo
k6Fe/uefiUIiJNNV1w3y65gBSoK1lfAKKpllkyjuz2oKPyZ3AiUoLfQT2YAA9cHsAdl//aM8QDsh
QyJILl602sAjXL8/Bagb957vfVRufcpizTCGeNRYbTsU5F2OTAJYciOdrX717KmDBHwExr35B6kb
meUrCpMMVkRWvs++Fbr9hteBhqcrS2MAIVSeqxOgNREqtXwECigiyr4H558NFofDBOEhNs6G9giP
T1bHv2BQ7flKNRLdtKDCFtrUsgKQZ+pr+SflVjtIcFuKOiVl7VcZmQxRqhNWsGFBjpbjLbHeXBQz
K5NgZfm/vjUIZyVtrQBrFhY98dO/R27nrwd9safssV227dfsUy7uho4yZaf+KRKAd6rbGmAGzrc1
rglGqvPTkVcHoarFfjiFQzULNK5+X5ylq5iGM9rMNINU+Q2NXx5TexLUPrbW4ZhoL5Nw9/7Cb/92
F+c/R24U+uywxMJFQJKPN7J/usAMaTYdGURMFnlcGE0GB7VNulfK6qrf906BDbzecU8MMm3rLDmv
qJ0wbXVv9cyTMnIpDnDRRi4IH3rWqFtaAMwLvENSAdn9i1PJfbJ3pgCPND5s1L/iconm+6Uvmy5a
GMf9+QhjKliw69tCJAYdV4fW12d14Ugyks1tvwvSIi/9YBMAxnqeguIK+CUIx+05mG0vYH/DAOrJ
7HFqEx0P3IJP7AAZPBAfq2U+l90sTg+NKem8U647oaU1TbssRvHRd6tij7L14HeaS7zFo+ZTeyGX
GaH9vyMJ+X9cXniew0hJils5Q8bvSRLshCfl9+zASrr8MjEOS0b29ka8ZJTehDeigmLLHvenDyYJ
2BYL/Dvj1HioGsHJ7nKvENPG5DepO2jOqQn4uRnQibqcyy3tN9wW+aC8v+l9+s3HBoPYQXfSWRAC
cWCFmOmEEmpxx7+djpKTntTRt23ykV85p6hiv8IE0hOopFsnHLMACbfbJMyzflakv1ekV7fY1gvT
mqe58DtgvCeo5CiNKGPrMwk9DG3E+8pXkIsOEC4PLZWcihcpuNhJQzmCiMBNDwMmT//f0KXWj9jL
DqyTY4LOEr/TobFxM43qioIN1CbhD4ie6jTUsxCPnvyhFf+pYkpD8IJRds8mCcKGZhJo26YnD5qq
sowvyAD1sjlfB8tgH3iAxDxx+vAjMev9cu2ILmr4SAlE7F4JLQmYOWGAkztBUo9CRXD5OKiSCN6W
DxK922JFfqDpn7ZYNAaWW49Oh1b2LuExTcIUZ394mhpGzfua7BrBsL98zSp1qr3mMa6UamY/W9UZ
CkSvN+vRXWyr7Nt1D/hFotaer2oYpjNVh/xjJAQNfUJV+qkq9ganzlYAooEGERtvN5Np4wGWo0zY
RFLLOYABla/VnpVqNu3PSmLKkFTMTHIpx52GEfpc5nU+TDvI/bPojFrctTe2fBwGtOHPborT0Rmq
8KMgArvbDgTYUBCr1YKnXTOqxIC98/yLyEZHLsYfA7cr73mQlhsO02RVzzODuFanjCX9s1wHTtEG
sJvytLxGW1u7obBC3wv70ReTxbJUbwHDiSZ+ro2y95BKiLDg5w2oqkWqElYqvFAZv38zhMhFizSj
u4bZGVNLeZ0a9BNLoELdUol1lT2HYNNHcF/STmcjSyuiELTdLKU57TCTcH0wZtOOO6YriiVMaE4C
hl127yd/37IUHHoVjs+vjvBfdBDIAoHRg0xEnBHOIwysEwWuiENBDjOOYRpgCf+iZbMYbhD5VBJ3
1a+oFjp0kM+zfS2sx4LoSHz07/8WcRAJESwyXBRBxfIBmEyji+gQhlkPDOljHtjOnx4Z011Ae05f
SWZPXaQYl4/TZ42hKwNqfkgDqb99kXdG8NZCMnp34uEHNH7TTGQQnxbzUSYP4wOGqxzX0EsgOJSM
2CbHl4sOB+D3upm9nXZy9uUdL1OyaJNgL3o/zoz5WvEgCz/5ALhvtZuRAmf/W3ZxA4oy7MCnHkUm
w+ONiY+TBT+D7MEjey7bYsrX3xmO5Vuir/VyOFbq2SX3ACyI419ZD/vuHpsTlKObrnk8H82G+Ljf
C5nzVqt3rnN2PlrcGE1Cj9vqrUOZMLdVzcdd2JBFZEK9l+g1NJngkTdbdwv1i6LGsHn0rloMdTdJ
ayr2Z/Gxx4CoH77EdVU291zQgCTHpAnJyopr7MHQZ2HErOfQbxZsqIT4StyykDN04AW0ODv3D3EK
w52syBN0bRA5iAVNv5XOeyH7FuFDKlXh40Wl8P0IK9e+RVNalEtFucq3+LjF8q1Roz7U7GciQQ+P
xYNzLSNhHivZ+u4WrEPVyMg+Byf4oAZqsOfNZDOi6SXURP3qiQ+a3UZjJCwN8QQe7C7QWy4+jLBt
BZ0LLMAz3hT9XAo6UcKc4uoL06qrUFkANDyLF5GKLHcSVlV8ub7mRy15LbL7EHgNvGNPVNP+FhTC
9BS4PeUxuTyccfqDiIdKcYXmHgJ0sD+O6EMMWp4s9uF1YX4oidVp3utXOKPFpJGp6mgXbN9sLnOA
ggHzwih0PIkWKcNHL2yBuq9xeu7SeT6Pt7+cvXKvIvgUvt3e8C2Xl16mp1gLj3GRE7GU9jZR5MlR
hQhYVhXSo0u50LtPcD2sbJxfosn3XUrdomfvGufiFBmpF//OGr85IMVbwlDbr/FgpC76STs4P7nb
NtAezQrxTxNZ78LGUOyaoTnlhDHTLQ5stOr6QuZIGExvFR8rInJEAj0BXUKUQXZ+o0EfdIYViHhh
5ROx2o1BsN2mNIyPii+P+FJZMZV7+KPgRKjqtCUW3cKmA+Zy0IyrYTfOfa4c3DqmtKhu3fdBiDjo
ubtrZ6f2+kfctzxc6HNTlk6qiy0/rpR7JFh9nadsger6YusKhIFAbLr7Mbcayd2tW8AH33sx6ycV
1ZhlTv25sP9A8Zo4BOLEyZD0C4IRgfSwZznmZig2998T3GuHtRTYME0xmQGU8y4mn0HU6Sf9Jxw/
II43CQk31nHYDoTlJ01/BmZWrCAnlpUywPRAdBayw5vwFGBekPcqJBteLrv5qlq5KVlyjpwyTUyh
v9qXD3wdfduSqtxvYHmyW0g2q4ioBF5X86mQ5rX9a4gISEBhozhR90t1wvMiefVVcsV6ROIlycoW
FPva7QOcP3ne9iSnyFOoHA7gWidj+quM+3lU7JZe/aCrewHO22hyDZn6mIYqZsVEFANB9V3uEEGB
hXyvRVHYoQ5eTEOat+f29xFghTrvHFYhuZwq5ZnWiDMB1An39y28/ftq2/2ggc6SBexq4IyyGubw
6z/5whbN6VTm4vhzUB4Mfm/KR3OwSnJbG3jcbGJzOc+1sRdfwAouBt0emvan/1Lj7FqeK3DG5HFO
6dHqiZzk76nBDTwwFGqhSpXM0uvtl/JcoIK09YVBuEeLscASZ9KRYAdo3f20ziASMyUA9GEluYqz
YrDArP5k9C6a8Zn4yrAXYbHxRexOej9D01wK33QxvW5YNnsDmiBWCWreZ7CAZeJUj1mWxAnb9lsw
ADwPFYJfYbq8Tbcpn2YR4UuifXSsfg0HSvb57ITWd9vpruuXojMHjr5npWzAMYFFl6gulX8K70KD
1U/elrq+Y9XkuJSBxxv+9sb901lKPoCV9F/h1q4BTuSUh9VAhllq+OSCMvsLLnysnay6dfULVlue
r6pY4vA8oLPclvreGaSM8Z8z/wfQUEkWWqO0sMImImcoPdAcFPn6kZpP7un4FGA2yQxeJvrcuqMY
SnD1y5sSbGbzChEtmAZMM8HvzbQtmK8Rk34xTsP75fYZo4fi8kpR5HjTdt6ghl6oqPH79jRXNKOF
x0vxcKBohD4R72fv8+xR6KC0slqzS4b0fj2H/l+4gT6aqE1hBn5cWPUDWgujEmdrRF64dDwh0aV5
jFLtjLtRRuAYZphYRYSiY5v2uAOoRosQm4/x6ZFe+PEooUTzavO9/VFGTzNLjOR+M1cxlLj6hc7e
qXfg7AwODenTKnoAj/zgr533MOtnqK1fJotcJwUSwx8R2pdc9FAmuETVVHjRYwqqzBB6omf9ldKa
S5wbo2Bk9NvkU3ax5ezIjpR/dBqXzqJw8Z6k4ffLOyDoQ1nFkLal5RZnyxemPxy/g+BpKO1w2eKz
Yzx9PDM5YHzFzwfMoSD16A1bA74isjJhSkKjbxhbBF7jUYCLuvcLUXLkp/il3qeUW8Szs/Gi6dwa
S3L0ngR10m95oUJyZILxOlKwkaEqRnkgo45mJVFahPI1O+DgMUJSNYS8JzrHuaYCRdSxxTPlKsZ/
bzDJNgQTTneeJ44N02HxZPbj/qpovJwNsu4kuROVfRFq8ADzLF3IsehuBprd3lDdxUa0dExkPY9i
kzjYAXwtlmZ2UhbE0LbhbHp2Q2Jz456FRXYxtkOiT8YXdd0JAjlnSNTf00YO9Wy7atz8XXEvJlYV
l7eYrLBPdy8bZW7PNd4ZAWlB2mTMOySnLmzF5ib273tiRvHkRu7DfI2xLhPgPpu/MQlyfTjGX4x4
ToGz8aqkm7i6lKYHA1ivtbHRqguh06/nEtlAVpCnSrsk0KPlcp5LaxHfkxCfyxCAK8s8g8/yhr6l
/44NE38set2hhlnYuOG5jiGvL5aWh54YdIe3fcns4X8fqB9j8Pc/T3YrxKWQTewPg+oSFLQ0tmbd
wAIZ7UBmU7+t7+NifUUd6j43k1G8f0zMFul5rgRyOCZsSGP6ltnrb2vZvrR+9kytS2l3oirnft5C
ygZ7LsiazyqdXTNif1noJJE0e3CQILz+vQdeKEYz7xZE5i6VLW1hKdJ3OpMpaX/mGwTMwXTKpxzB
Svuh4IcsC+5GzA9zLH53TUEEvCcBBTcLcKRujIl200hkt6C8xqBUXGfRIPTxZ6g+CyhKPDTf6bFH
PMb0K0L5lWwIbYaZGCPN/SfetZeHT1a2TjH2m7FaUnR0GgB4kRWezIsoPKpGBoXxL8rrNUsyTNlX
be/aWA2zAUpgouRJphYBSgZ4xWDMC7vo8s7grJF5gpZ4E8F7liNovu424hPfXR4XGtdSGC56uD2t
sgs7edkxn7ytExYpHdnFxwLLA+d35MSFfWcnxPQ+HUmemP8mTGtyUYi4YM/gRf9lYsRsHQvO/kq+
P+ALdl1VUbZ1nMtFLRvdM2eWj7cuJ6Va5POm5c6OO28PjPq3LO04eLNyGoItbM0o2kbZwA4IPhyl
bXfXWsS3cz/3yyUfiUjdKrOT6xSRWXHg4XqKnIdaICYagXyN1O0l2/zlMin8S3WSue7ZFfN2yMRP
VAAC7kA+j3pTTJA2cYAl/DMq7xOjwcJGywtwAiNd4Ao0Wa6sfgY5yHhTE1Ho3IHzJMPvWEtb8SJb
dnjZlwnWPPkqQyXOFJPRJWfiqBpbAQ8kJ6ZrzteUaTqp5/k85PmvV2mc9zAuOOxvTNuACxlv+dPy
YDMVDUeIIqqc0ujZTIrqb3cEkaYdTWcxvsm4+zB25AIN4ACNwJzk1StwHblPofjAXnYUYaSryzvu
IebvNjSWrXQ0RlL654EPP/edyiPeJspvmSGowX5hxCqNaMXtfyOCECc3pYqUEQ14Hb3o3dc6D5AH
WErdO8Mcyf9LNwcCyeHxnp/wUNnVBi+fDo3MnRqgT0uX5CCZtuhiBnp0d3bjoJHAQmB0l5LKSLQW
GWlHPGTSEhjdvowwM3b5xESaU1oMIQfn9S9AIu3c0JCHcnaDCn97BEaLwzSzkw8/fVlPqFup/RW9
eUnWbmBQa4Gys8Zy+jFiKwuyHajqIO+CorJN4XVtXLXWp+5sec4sfVd3w1WtbzGTKylFNSw6Ohjk
QP4DuoITH0lf0w9WoXF0haO3MK3Tyi33lGtOy1SH1WRFYcWU9frD2dgdjiXKp+e7mu+u+c5tY7s6
oeoLxUhStzqS31vPWhpm85oeRApB+eFDUGAxxmrzSOvZZJ60fH4gAiKHig5HhErkKf5YSobac8PU
M81NuG6n81e0bOP87PQH7tHo6mTNOBUCmMQKyGWfveY9F+u7lQfUUigsENDqHDKURVu+4h4O/NaI
MJDNq0rL2QPmVgigsZ++SgIy5ppmY3+hM6Y1uQ/wFO/mWwwkZrVIcIrSs9rGqXzpMd4EXGp3hxQs
P6nP/0ySx1xD8tlptBuz98zTBLAgBiesU5Fd8eHBabH4G8oX8LSta1GJHxtDcuD9XYB+G10G0UYI
jOTNgmCXeBGliMrtraIPDokkZuSGRUu8sOnycZhpCRSwgy/yc3Y3tzDJ84nwcQ9w24VCVfuY5uct
pjRYA53osyMWJZpSLLnB4QWMAp2TMcNbXHs3cdTPaHOeCo1MUsP1Gnifzwp2XQmEmGiYlf6AkCoF
3NA4s6PML1P+uQVW7zjw2tOc5Q9ZIzux0BDuRdk8LfPh+GtEjkPijezpd4BIFsla9xXHjqUei12h
Q2B2fxVzp1khqeAe/e2qci81BIoCS2Eibz0vxMFd8qKVcyrGble4ISxrY27rkOCS9qh2ioduh/u/
6oXn4ya+ifrWf7sk210DuIXbKDqo9riv16HovK+t8LLkLICa4KbKmnTTNGr7Nqlm5ALNaFw0Bslb
22rpptYSuCnLM+bxBCaovPDXTzlhouYyonEzm5NQ5kEqcFrayqE/0XgVO+phZQ2L0t4Fr/0JNzip
rfP/GqMuts4th3jgqx/O/xVwnF4oJlkAUYS1hRCA3LqpBUVijLJFWmJm3AS1i0zS9U8LW6rtSMx2
BykrN0AZD315ZcAGiqIJG0k+3EHVHQF+Fb3ULart0ZyAqzeuGXpvIuvGMWY37GtE1Sb4t5WZal9T
7QDR/J8o0kcuk8bhaQ8MF5SPnaGrENREsPnRzlcVlSGHKrFwXV8Priu7sQTuXcndsekNIkuqnTlt
f3FCcheWNSOilmkEIY7xRc7VN0Jrkvw0fwiMCQfayXh9EkD6zkI9C5dCiTxwPR0d9tlkQDsh3RRr
nfU/F8hP16J/uuyyV5ftJ5ydr75XX1LyP93DUVZ8PvBbooI2rv1tQcL5Hh6F3nJyu4q6wRHuletf
mBj0eZN5q8W2NuIoMvtPiuGxHNmvXETiXx9AGffwJk83yVyL7oUH8UizsAYXijn9enAnnZ/WG81w
3uJ3fGs7C/1eCQrh8Dst6EhCBpNgcgWm/ZibL0U4Zx3+vHMfuJaTXJG7UK0p5zmu4YVhpKREX0hF
dfFnUeWt7NecfRK1vcJCFSwHGPNKQj/9mENyWFQTvGwK1h5OTO/HPO6UQQtI3VcSE+ajXRvW+hwx
CGDLkPQVHo5JMwulkqjdkvIw/yEHpk7hy/XZeZZREz7SXZc2vTx5LP2zY3xfrPiCKNntBPTwWqeK
kvnhlSpZLfcUIvngTu4tPOl4GKOTdGRFPvBMrPvP7zCip3zJTeRc8WtAU4cLQBgIcbjpx/1Pf6RL
utuKjwwL45PwyaEcF0nQNe8srcT7Ow7ZUP7kkaQ7/0xGd8578FEFFBEbfBqRMzHV9RJvLWnko1ww
WVdgw2qNT5YG+mYHeCoyJhMaK4xSnBKSxocPgldFyLgGvE3D/MmOkNSdaTZPSBf9qlkz3SDEuQGL
rDMQK7c3AMsH5v78rlxd2AxJIgWX4NzNuVY+g3VvfbUfXdBqJe8cusq+l1IWoEq7fq94m6xUZ4qa
4JFixO6SSKiXRChmA/gFowcEeC5AKbxMt6CM+NIKoPfCCmaJ5qVJ0w4Y3QwVLELtN8yImoQQTHqH
3d6qJ2YB7eTVv4T/HeZ1QecA2+3+1J5oQnKb9Zs+HF6I3Bl4rgNNU5Dd/kYdi4rr6XSnYyISbktW
59cJ91ofQ1B26p1phx7VdovBiqQJm63y5sbFWaOrlFtYTCEfmLyvd4EyIY25FUG9etKSTIbc2Ifo
D+OSZZLehdtgutkCM4TTMrYJfKXahh8Q9lPDJmGXf4zhG6cHdmXr0lAq4EiJQPUbHpr2xBnZfgH7
ZmpN5daeJDeQiKCBxvEl4x/D4rmU8MMxpY/vo5af+vDm7rnMP0+uOgGQR+aTYxO11TfjzSn77CdW
Iu1dmoz7JVKZBo2Z1c4vTxrEG57LhGTl74cx8aqYBu+zy6sK4kLOEC3N58uO68JAb0P+tlDLuk3y
AOr0eqwuE7LI8NrEnl4e6JLbsV3aSmyC4rphWDR+RgRPvX+UiJDS32WgjcipcOiLmqc9u4CdibHE
COAeGDHkzIzAIpZMcAiLAa0ax5tYQ3WfVb1L/8GDyXzj6XgBn8cpb5cwL/PM5MwrEW1fb7haUHVN
lZquZUpeCAtdI495m2DtBCSOiIWn3ByIMkRL3YHgUJCjm+cF4QSQAzUVk4m2GshzrxXj3Gr8EUsy
htvPVk8g2yAgP9cK2XDt3A33Waym8EqeLIcuwIXhkvTuRnvvT7B43+83PlAPP3vDqwfrwqT3Ueho
me7sFltxaopXQVScUYPZ7jbKCwi2wDzUwLY5gY9v96Qp5aYpG8qdJPd8sKId0RkeiPoDzg1SvpjC
HZYDEjK3Ososmn7KJxSqHHK/cYPXXrLNl//+Yg7rCmSE0w+nTQQvpxVXL0dUnnGBShHoLym6e6CP
4b1z2O6dJ4NBaQ7Y8IDPkscdWxUJ3FYdEekdhNGy/8p/e04jxhnSfLL5gkDjWJjm3NB0IIH1CL9w
EJhVzYO1O+Y1so5POagoo8oca4qDqnhO8uVNiQ/Spu9XektzMedUN7Xtzz+oK4ldlftNzmEh8PN7
V9MsynD+4y1HKTxI7UFKvg2pIaaqRW0Xtf7vAWobXoHDoKBEmD/39ZYRf+Ho7OpxFllBtqGSbzZn
JqB1IPTK8hd/6/GspWWGDp2UsW1Rd6t1tbKYPF4LSUtLyDGhPAFVUvGxNdQcZxptzfJGqIKQTO/9
zK9W1981GVqpbvmEqwp8qc5FJxmnavlYF7o3k7Th6x/4YYGpJLTqaz/gaNyTkSpr7UFTxpoHXEVh
wDyd4580K1/RoUU3wU9GG7MqPsTCOk8Ah/E9sOlTqMGzxXB1SbIqs3/0v/SV7BO+/3Jngat/BGj8
n1JJELchwv8ay956E2UOLE3fOAeJVTAJUrJ28IMG3Y6qc9XSI1DgUSxqPtOjKmKNxdqYcEQqUnJn
N/0XLQhQCgMbr+qJ55VtJmGHxdgluCgLq5cp+UbQtrXXoDj6ff9kxR7ECJDeEWlmGqUJG7YjrjKQ
Xv37zCImTSoM6aEwpQJVXzageRfEITKMits+s7fOh2sFGQxnfXqEZ4ev/WIpzquiKtoGiomLSh0x
haZyLH1fmc1g+xtiyWCyNmMmY3NQ5X44P9WGZZFUuFwbBJ3rXYfDeCqr9SwfXctCHpjMPT6nefdl
sRfkcglv0Zp1XY7gDeNdfVfv+tH0BvO9X4C6Fg5nzVCCzukuWAL9Xc6KIP22XK+f6T7RETZBhMoY
HIK2q2s+Fr63sV2PU9MEbeO1w2pbg9Xh8RBMqP9kvJbYENGhWhHGxOfQahaqlrZIgEpOiyr9Bfes
Td1qRsOlCkGQyTYGrdRsCH6HK5+Pa+iC26sXmbsIclIe1Ycis928zoiyMQpez6kpnKwe11lSoVR0
EkS4IsIllcZtuCQYGpsdMh4up+slub5vLqHM6Z2kL4Fpodf6Olh+4LYC9it0X/K56ds914u7+mhl
mjrywn3RmExDuzzR5QdR9pog7nisj5i9u7xn7aj5xxn8zRTxJutdikIM/hbJ+8sRNJKGYLKW2oHx
manGEc9WyRF7xurwhPguhKzrtfpgSnHgkkYTIaIp4GF9ttPBX8By6fNkoKS8fu924WQd2NlFVrb1
Hdl1x/LhRRa7aJXs7hEDZ1ahIsz6SJH+YAf9oEDyfdQS7c2NMRnbcVTUEwUG1/jlusApZeqTelbT
Js2O8mWgShibp6/HLlAUeQLFAM3uLU0+3QbwJl2EyK8pjRjEP/urND5yJi5iu11972L3vE9TNQzL
0+E5GIRdDgncPi1TbjaFs38vANOSilYz2ytUa7Co+jVtNbNODi2udesmbWDosCYpxJjrA+D0nVM4
LJyOv5Wr2OR0t1puqBb5zFMavfKvyUDji2rkdgvMoHUlNkGvPyqmTNwNjLlvWXGrgBQ1P0YF04k6
0/43b0OFLXouCbmTtJEIGLOI/vetn+gkkhBjPvqDMHJkaJFEL9fm38lcZq9hA5PN1N5MITpKgiPF
c6cUXNoJy3cLX+cZphEeQlOo2wi+zbIP+JwBMWGiLke9fizLCoEX0VhFy8rlLAGKAUqCWUlUikdf
Uy62c68fM4vPxSdPhPpKJhI0mtTE+HlVFryLFvbFQbhOVmCncpL6XFpk8xdlA0l5/S1i1XqVAd2Q
fbdujIY+6IhLSzQS+qaH53cX11MRgyXkKJdoqlsr76arSZWMRdNZYO5Y0kMwuuM6d++48IIf4erC
7w/KlqtAwHJXVuloHHgJ6Q7/5h2KZgSL9O9YspoAnR8tJdGzDjoRaj9gE9H5vfJg5pCVvy3Von3d
BxdLNkoxMCwjfCn+pcJL4/7reXh1ZphD8xLqmoGcmJ+dSDLszq/HodRoxcwe3oGUEodwgw2q8Mf5
oyxc+whvsvb6DTc92LQ3RrlgFRi8/4u7jGGYuVAFbdwJifKreC/M5DhL7ElQGm+dMSJELOB5sphF
J+MggHtfXOYZUQa9YXwbDp5STMCUCP/RnI2pG8htbZIreuPDnzs86ZL0rXCqs2SexySzHH9wmdg8
CELkXo0vvGFqPATE7gWTU7oufRIUDC4qKHH6zmr6+/WH2Kbx31N2OXfEkgasQK6gUi3crVGJrH3V
+x/xYA8UjBdy7I7540zTXeuxH+aeABJ1OfQw/e+pChV5+4fgnkWt9FVRGNP1953g0VjgqNS2E8Tc
5xl3UrHMxA9pcEKL+Bgq2xwB+6ar961GvYuVUcJl5qOvBdUyqeM074pPbSO+HD5OaDZhLTHp8qBN
ZRT3YZ9iJ9HrDfUA8bODE5rH3wSTX6VvmwjZn3ba5kX85PpfxQKomPg0yinEAAeOEBvZnYpGECFc
gXfU30gHAT20ntGUvxb1MkxBwyMPfCp+WTYEWM4BEeT4FU+8y4NPetU/8o4zwYAoydQBJ7wT+Jk8
IQvz+SkTpLTxFn+NQ7v+hemEnl7HbiTTiYZ0Y3jnpk0+KvuKXHEgYCf1r7dg/lriNlhXjlwdAemS
vaM8BAlsxI9u82pdsfQtFf8fm5IMIPtkkN+FE+t1u1nN7IcYmrHZMfEHNreEJ+qKwRJr/Xc4c44r
ZsY4RlNu/iiJgEgld3HcluG3Cb/J3CuoKk94yoXzmKigRe8ECW1TFOBK+KqlccdAQDfAR1hxnaAo
LSGt4Es6uy+0VhqILA/glq8E9SdNPGKyXt/gIaGA3u62l5+piBBD+xrc2+hMu+tO2rAapI7/nSbk
2mQu5rDt7jLrPlPOO+9mzH1SBRcFA+aDFxhY36btDbeF31/BsLra9Qrbqt8lu2FkhA39mZBF7kLg
3PoLuLpBLHLQrR2fcv3g8ctP4RVzNpTxdcaJzbYGvVCoIpZqjnjUxN493byHNTd2xphEEkaIC2sW
haRkIWv9naDIAxEsWe6N6y0vULzi0OBTjYWxrHuUgDJ2BwlL8XWDj07Nfp7RQS/yIbb7GF4WBQGF
Bl0KwzWntT66VVe7VJQPiRJKErkC/artiKzHt2jle+P7djibiU5b+GbJj9VauV8vow/7K3WuWUvY
JlGgqc20pAut/mJYP7YS1/oVNm4a+dmDJKkX1Zmfk+lecPG85mvaN/NoVKm1yj+sD/yZieB22cW1
uCtxEPaYkRiIv8O7pJN3ufktXZN6nU4keSCFHxbliN+d1ljJ8HZ3eOn2iv12ESfN/ZK2uNBiCUNr
b0flSw/1CPpnG/qbuSxurTLY3yfFWVzBh/sJJ3PjdD4hRqbjNUVC14MqZsJJAyDnsGOzoi8v3tQD
VA+6vshlbL+eHg3Tbyszbchh4ZwQ+cI/9oaJqhhrgMgaUOpoERUTH8rjj/UyNNDjV23Bv3JDDPLw
OQLRoXvNfNHyltWwaHzlZSTVJ003adRemSVXuPy21J0hXdcV2xJtkRf9SAJKAyMcZe/HJ7N3wGw/
20NZ3lezuySKpuX/kS8Ub1C23TSkQ/+j0BnqC7lqL7iZbLShIYk8jkVEOdbdyq0qdomsyyROowEA
EmQ+gum1gE77inyREaBYuPFh5eKzyq4Z/N7vDZC/MMjLkZGftfoUVgOZ4AVWc8LxHCYjciuu/VGc
W6aw3xssN0EvawT1CWWYzJDUMNxmlJrtEVCX+JWj+sOLcuL8lzO3d81KWZxAxIAiGP7B7wD9iXmI
SNr+NkR7SES6o75GoMx+Zo71OgHEN1LnsrTwiyif8P3YlaM455SLYLMXCYTukbGi0Q6AIpF3TZ4M
TSMZHjBRKIVJQV0K/N7HAxGceZCa7OGlpwiYyHhe1nZfqKAJQAFsaVGNYHZypnle3xj6ogEF6paW
g5Q/8j6w8tyNpKBbIPUKSC7byncMNnjW2l7yu6LR1R4BO6uZJwatEoSDUAWqSk4fQVXyadKh+WmN
dIgXJzFxzWDb4jo/xTtNzjc5MwbUuMXtDQetgDxC9Yvh4rV8H8hKdk1G65ioJlE6uWrM9XIUZBbt
fEsc0FEFXUL374YXlywAKDH5TXRvS8eJG9kXnkBs/ixRhuPCct4NtBvpNA6QUUuWJiRcUKh4WHL1
QUuNxSH2HnSzWkMPjyJUoNkH5Xxxcj/cfSiSsQYEyJcQZk77Js3I2n3upqW5keVAe9HSmDhxzci4
5kwf/6vFz3jmIbhaeELJRIfBKXkjypN/jCMpYpCc4VjHbIn4NTZkpAFaRO0SgDAhXq2Y3mZG41Ix
eqmxgpn+HZsmDUVYgR42EF6KdGxRA7Bz6LjMfj/7Hvp9was+thqDlP6KeJaW4YV/AlVLKmKEtk9I
rvxTEIOj7UQfZq2x7zmPGHZ/rmdEqHhvno5oAj92YVttxZlCfUK7GLgcuOjiveuU2l6fMoxQLQ1o
o7DkaZOwhROJEkk8HEy1MD84oekgtgaTpSUgacXHQKRl/e90vJ3GBQoJX2PkpKdiK8OzpIozuySO
5upn7s5kHVv2mjqCPMuz2Qvrn0A2ogGiIS2ChiBX+JWElPzW4AfEELjB4DaxPlFsVEU04rfEFvsj
tS5L2i7uUUN47X0QFCUzmuA5aHYSZnxnMyO7pt/MS7T0H9DTDcw6M+Y0e8B6KnkB3V2z9tzkbwbM
fih0ZAFlCOqQyBBnWx76phNhhX7KH/+abmiZrBpWsoPHDg+ItTjvYPfxGqXxRtDdnDm2BNN92+am
C/K7B7zBn6xZDzJyM5Bj/7cAU+2/s6oKN3kpbmHXEOOhmrrfvI9/Q0rmFjSSwz4ZwbPz8JMjuUA7
0boI19fFtho0pfgI484+Y6UwOjBU6oS6iU+RdwD3so81HuPNCwBq8oMZ8tXX4FWcNu5wpH2ArQnJ
RtVmpIb+ZepEpRSuxYLxtXflgxwBuf/ZuTsQVrh4VRzDEZVCd8wjFVH1SHsHlBcD94m9e3ap+Ki6
VfclAD+6QJKOlz8pQYWfCJ1rQnbeBWWbW17CzsH+BCLqBpPczrrKE8PPLKH512eqkbDF+oCsV0OW
Hyf9WqWsHjPIbUNyN1vMHdFtODBwlw0wDb6RnxNCthwf8QnAvf3YkUSW0adOpc9uPxnmTdSbQs73
6Xz0kihjj4wgxRUJXM4FiIcopiy0Gu2Pfef+ewCT794VgBOec3vbB3427hSTV70wixSJO2h1uTGr
RgaftKfMqsKv66UrgJkfIfCUlVaM/F74Vld4Mrfy5AeFuJV/LW6B/hHGjGqkDeIuZVRWWyDlH2ed
EEScps/FJ1QKnQLMZxwzICsb1BW1PuJ1B0nlgbbtrIb5R1sXVhm1YOW0sAixoOLkFOl83THMl5lb
hnbq+Tm7eFiyME0C8mj+XQ3mN9js2hT/xqlH2i+NRwpRpSt8FAClHJ4qvx2IVidaxWa0C1LzaEGN
R6OlCbUTDm7sKATuCDu6xLLOKZgowaIjFZcDETsu9o0zuaJczQB+8utXpJ5a9ytwYJIvEmyXqzUd
49FW/Onc4jgD8aJ3AyLb6usJNbwgPTYy1qrh2r5RwSXkB2Zsuo2cJ8YFTYjsMM83YPC7Bn3J15oX
UcdJDzZjZCoRr2iHT8M1Na6oBTWZMYiw0iJb7lRhF+LePcE8f12966MKKJNWh5PYQ1smAktpXdXu
+i11RRV0SUNjHssdt4CXFbanMrXiff1mlYlOdociN/wy4TzhG0QDoNAS3S5FxWzB2s0qlBMkeoY8
yWSK8kTSU3n8ME6/F+Hsxibpfq++C3AeLq6RgkSmcqvIKpAgVzKgsU58VfAIzup72OPXh+0QT70u
0p+hYz8aXqBiv84HQDC3hg4LZotO9VRzpow6cqen9py3kz9+oxhamTSFx5IYcbzt8AfbBy0EodO/
fKJ6hDaouNE+nekcOI5Ze+K446IyTAgcvEf9Bt4Ea7isrHL4dasC8ffySuiWQ2SCcRcspyFrn91V
TOk46FXvV/dRbP36uV2UziN8NSk9QbG/Xrz1ZowpeRzt/HSTOZd+DGOn2ZN4KlZ3hsG+oQ05W1d0
ySg6HCmzbmS6Ho5q+H59KVJs6CF+K8uTCIWhesAGlXi/vrkYhXc5Uw1ZcCsNaFaeRlOiV/cyPELS
+9R3u7ej77ZEc1L6RLybCX1hopx3zoM6SGCdpLaEu5X7lT36hSAWSIYWScs9RSTmjMv8il5d9U57
tk+CKoXGAplIPZhUmSCoUDbdZXmYXJYHKs2YxP4ezPHuZ8wFqr3AbJdDj2hHIR4KxEFsBsX+2dHy
BHdgDXNnu2Kd6HLwjUKJxNbFSvC9BnwvVwXigoMHIUEFzSogaVxKWuEEgQ3idwfPyhbSB30CxNNC
jysazl88m46bOFTsPrnqTdEapZ4SzxWInBCC0damythL97hFET2gnBNxkq+8whmXXWfgx5WVbyJQ
mG2OYFbsvafhiX5RVjlHGVGTQnn3DK/x/xsGMn1tH0AcNRQ72RNQzIIUNdZ9NkazNixKEaTtn+V+
fc4L+YBhQccNI3bJGN7i4XkoX18X0k4/cgGd4ECbRkI60dQ71YJOwDHxyd6H50qFu/cE4XqLyqoH
0QYamd7Fk9OPSXiUfU0TirhXwmwBmUsOyqKQE3meal97jmg2ju0dW7UBVsK0o9jPNA040pCat8yH
c2Z7N2QdsIfx4mudalGtMPtVKykoTU5FQ7P2n5U+mRitq8hovI53NXVzN47B7uvQj+3B9sbjVXA8
5VJvolerivq0xfdHP+cHZgkYwP8nkbQQrhRyk4n0UaQ6QudMvCEWjsRVbS3x7YztIc7hc+Mh1YfV
YW1hmHnXefxsPpLif8LmiZ95m+Uep45Ly3dY1Pdq0PDRo4Uy3SwQyuk4sg5rv1TvolSeUVjy2S7q
t2XgA+mk5KprVej12JPmKzOgQYCXpOTXXKlwvxnnD0V3NE9EMGx9zd4h6GF5tvxfJzGFhqoJ85If
I69MoZatd4b2ThoIEziEy7hWL/0VW4QRuR0SGcV+Ey41xrgFhKgpi/GIJ0dcYmBFDjNGP819Xb5C
VRbDLUVr8JVweVM3oTocu3sWoDqfZdlWvQ89kyHgu3Q2McHwQvYJGpwiTrsohxP0YGixB39qEPxj
wUFHhm1TkZpSUjrzURpxMOkaTPGdcZqtsyNGhn/xPtCkYIHSk66y2KuKLswek56G0WSxJVk9eX7j
Fl3BlCTF0E3Ps0ga3tYmgk3BH5J+9JzkSD9IkRn8ddfIi0PDO3upX4/5Lln6NpvFy0iLwfJlVwrV
WnuuypPQ52VdgpzGxVONHv0ix+K1YdD+LID90EA6VLRkGMIO1S2W6zHTefaKP/L3yOH80nDRHBjV
S7L5gfu3RBAKIhS0y1gBVKdLMLOxK7qUT4azV7DHE4AO3NgonI7I+4E1hn8ObmQLrg/YGGos1KeM
q1RAiCcC5N37MA/zHK2OVnt9azuvREuA7ZiKv7dgFEe+Iih+1YGpsMf/hF0PrCo9LSgV/tLrGMlX
zlo5+pLZ5vDCFhwFTdKpIPYqo6swuX238neYBWyQK9gzlOOYvl3nxHkUkNW0He2jW1e+L7V0qNzA
eq+rlgVDl1Ft8a9a+pZEYfK1debQXKR00FMCJJGfsJMO9jPHJaqXl9r/XC8KvZiUBMUXTW4Xhcwg
Rbxx/qBjXE2uYrGVwMyCFWizdYJoS9DD47cYElWgUqY/8NAjrQlIIaFYhoObYYmwyW9coRtJmKst
zVyRoyW8SePB5Z/7GQTPVxsNTnv2YkLtGXVydh7Hj2OYf23om5ZZWKoaPTU/nA9Q3+JZ4PK6S8uE
tIlIevsx757XMCewV/gwbpSej5Mhp1BEP/TbPTCys0jSiuGvDhTomS86q68MbjcbwCuWGcF46p4t
kQ5TN2fsltv8Vh5E6vJNCArLg2S5PGbdZ8PX9cQN6/Jrpc6rj9e7YoRiRtLKRBFwhXliDdtHatib
nEnmqIqXlJ/uhrVv5pnmq/wvMnfSgIZJly/x0iPh9cJeYKXwCG2hfq+HFP9eUlwRlbuFEBlohNqI
Oilkv2lV3JWqacPEn3I3NrUni5pCUMEy+Z04BiWt1JrChbUD+356j/pISZTTYLmgdl61cDmZqdjq
rcDuRm+g7VjOqQKnmAVzYelkq+a4xZdk4UlqS9LnYHgQsdLoiKaYOqpTkH6gQKA8550BF6tn+UJr
7JTH3vUk16HHhWtMufKYFDJPlcDKA5aj8h/ssatERCfC/cShlqaYM60NnrcKjNzd1DCa9yV47LZt
makJdBxTBDZIwgnmMThi/CLZE+dYgdm38nHj/gPKE1W+YQS2Rf2F48MTuSQgBB5B/kuo2fkhqxdc
WVk8L+ggiW7zr5L0DROtAHpDvs9PeOJCJSvL7nF1hJk3kqNTfdaMdVzEQOm2+ZOyCTgjqVoBvTFL
nxk14GwdutVMDEQuf4Pg3qgB8F+i0G75QcCjAadyIYRVZsMwxBSycCUy172gOHpqAJzOFVvv850E
iDbfViLnLJaTtO+GP4Q9BZo2l5eBuaxTrvLxJEarNcKAlDYz9+lL8fLOM9eXhMc4eiFvMjqJzGUT
cuXjIiHwWerUuWK7Weym3DcW1tS6VKp+2GPbHRv+8IGPirDb90b1cyDKMiXph7Rf1FQ5DF5NXkwq
MyTR1EDzcpLrZQ3ieQK/G/BCZHAutD5EWok84NegOWgzs8jqNjuMwMpSTzXe+Le9Kozb4wGdmuWA
aXL+Zyf0PDcdPix0SVhKhSwU1VVSiE9CEPCRcHmrZ+EBvG2/JRMaV9sriceisN12PS7HZdJiVVHD
nTShnF5UVkp4vinGLciRSGfGjYrJRq8pQiMn743TQD7ZKtl8bj0mwNqEwAYJUGHHPfPj9dGE8ZFG
2u2dUlYY+9jvON3kDjQTuM+3o8WRHUtlzTP+U0B9f63uHVHurumPpy2IHsLxQsIzlYmn8hVzApA4
EVD+BHG4FXQqSRnb6txwY66aZ1Tj38NmttZ43YzMXz2F+WSnp0ynbaAKM0NPNxqDvZ6qQfwjpyri
OZE52S8SEmfJqf2hqXW38JS81swdOXVKsE6IzcBm/sRMDQmoKRikreo74QTdVT/OAiFvryQJhdLr
ZOkPYtWQifStStnqBn3+eqeZUrqEb+qDhMo6tqyy+npNRcqaZDZzsNcZoxNrURTZwp9VrQ/zsKKa
LENMTEj2PKzIMC4OnNEUT/VxB6nyKhV9R1WfP/8pKl2TsDkYaw6GPPIgZIhOTQEe119MANF6H2oX
bGf/0wDp3XFUcSDTqGRljrS9+lTrLZYTKtm+44xbBaxp5+lpIokoN37VN/n0EBV0fYB1uf3ItcCx
DUfwXoebYhJhn/pIxM7fLWFlEh2814iqw3MfgCbrJII0cH72ddZE8YPr14DbdK+Xs9XqhrvEvM4n
EDUHV5BTH6DhG3UF3E1Peq7zV8Rmwt6Hd916xMvSIjWGoXs5uOhvgG2lEUAcNL7gTQLP/aD4p8Xm
GCgVJR7ZLiZpoo/x65ttnavJ45FAQBxx8JVrI3Ko1cJTYdzXS8acQJMY6NX90DsmStXS7lTzJ+se
Bw+miBCgZOey7bq/t8RQ+U69h8HCdu44hti9JC0waKx24Y1EZiP1xN7X9bNR7Fe7caXymXCfExqo
E2CA2UW8kc79agEtjQus6Iw1EAlArdLXoVSfloTijxwJq91Ja6Gnffz1rMXpz3xGrG4PgCdBf1Rz
+vTFuaHDP10APXdwgo4IyC6pCXWQH2M3EfEcXU5rp9wTCza+AckL7ISAIwWo9RwvWtxgxEiR/PV5
bN0pwd624Rhh0sNSp0qdy1XUK/Dh4WeyCy1BQ1AMJOzlnv8c697ltGa4TVWwHjiehNDVb+oIY2bN
65XdX398VSxDQa57MQjtIflMq9fOZxDeSfpJjwIRjIEHYYtG64Zq2MIiB8zuhdnUx5ar+RJJZzgK
xITYrcBEbanoREg2+4CkXBvf2ksOXn7FVON/8yr45dlV6WwyyS+vspvMSm+e6MjOTSHQtQ2KoS0/
te/tlNLAixVGJ9hLVVRN4L/Y6LWe/N5c+/GMLeW4eCZSQ7tYMWbJYXeeypj49Uof32BfqHo0HSDm
7e9+fvgZVtB4XWSr+slX4vo2RxMIDkh2N0kalKvrC9VHhGKdAVAJlIM9UgaRBLk7sGOQdlG9vPV5
jT1eC+xeBmTLIY+hlWpaFrTsDpqbok4Sx9ePQdTOEpA6clK02fy+B5OMAj2qq3zNiPVFZpqHblKr
D5gHMB9LOaA4PLoUge8sOAfJR/y/qql+2gLyav2e84ih4tRQ32WIaBYmwkM1Rgk3kJzrVCivDK3p
+IVyVchKm1Dx1QD3CNFL66dS68DGSf385VVrHzpbNLk35mNukM7pNZcL6jFoazL5j3CHEo2vNdll
W4uItOqVGwqMc+6eLzFk4XH+Ax4WvmJi0KVKOryiLYIyczFGR6F/ovGwmyBazeU9lce4LQVsxDhl
JrCd2SB/cRO2TJ1xANTdVY2o9I7wr6apzXf3iQZpjChWqPL/zub0CfDd3pq+lQTej5ERa2xxyjtR
JjWmlQbFxSzgaKnSqRZZN5qAy8cwGhgmt+X+t0NogWexcMQYDL/PRbR9hgUKK6nLOAzK+60GVPQq
uJwiMRqwseA9PN6ZmAgBgcUhD9DhCRDebPp8uP9+5M7uDgH7+A99uOJoxzfRxuGEmXDhF6m/gWCB
fWyKNdxJqaNixIpIS3L/00pt2IRdt38v7cW/10mWUZ3YkPM0pz12353l1RaQcX0eI6VCcM5OLKPY
qETajMfXzKFb94P/ZZi8n7s/EcHQfoijSgjnRuAFU/9tiEf+2q2mJSVyVHinO7Uq02J0cqrkP2YJ
XTLJ2CZVIkb7Eigrt7MvOuY6TKK664M6drobit7UsBOtJT74qnCm/OVS1G4susV2Rx9jPsZwJFke
GyXkNyCDEcMay4r+IlCLmb8rSgvSQOL/FIF2BTSDx1wG8J4Mi57pxnyMu6XUaa0OfVeB0WkziSXz
L2wG0KoO394CZ3MFwdOC8uLYoRa7u7kzVSk6YpBeGF05Dd/DdAmMueRzDNtBfEjvYVewChrQ5jm2
IXZBRGkLqORcjt9r2iGnofB7OpXqZF5wWfsM49qBvDlGJU1qPaG9X4ZFKmO+wk2kYgHSxionefnM
ySm2HgRIDdJTxTr0ycPdAROEGkvvlsIUoextMeds4Zu5SaYuwm4X78CmNItiHLVpjYRiCjei4gIv
Xb8Olp8fxsNsvyfBlB2hTmt8UVAkctY/Nlu2hkKjs1zfzHO7IDqhEGPLzLI5bVrcIxikBocnMtdN
R5dz0oEqgY2HUeY7fsBIW4RZJFcWwg8gr83FjGpReIAeKF2bLgsmqqfqeKfOrmelyXFGc6FlDZ6o
GbY8C+Ixm9IhnpVKGzcb1c1MzDQi1faVzJt+bzBBcvSABxfC1F8MlZs0g4pVChWmqAEl9V3ekmQx
UDFdi8JRVEdvwMwtFvPlTM4+ftzHJgRiCchPmhmRGgYwkhjIlNPDXCf/9oyr9w2qz+3Ux0CUKRzQ
sUWfV3kILUIZMZxFbcfLeaBEInuDCwV8lrLZHn3cEEwWPO0GLWHkbjLxzmtbdKkvl+zaRVZ7K65c
+p7wXF+1nCZFDJ8O+qbn1ndeWAQTX1qUypQ+W2WFdTPR7GZqptjQxjT8AqxYUfLr6iHSMuubbC2t
QLBbB4PEbGyxtEG7cyaGK+OdmRhkXzrco8gx0cqKjZ61gc4cyRz+wg4Mk6PE6x3LMRxwDqh7eM3i
6aSXK0hlwA1lV9p9VpnHJFxBe3ZrnjfA2iny+Xr9ggqvLaI0fNhQEU1KH0TBXMGE3ENE70h6BFX7
pWpySzeSNjdelX7H14DwKlgi3fRKRS2+wsdKB+nBK3z3KMTHcFNGrHzRGpHiPphpBBPulkupvZw3
GTOfag/nfVjaM6qRy+rzV+qTt+LM5IZPoFJQ9GjZeO48SOvmeNtuHlpTkv8VQCZm94Qqko6utjzt
k2A2weHdxzKy87vP8vK150H2aZiivXNbyUxN/XfKbcOjTXRRGEUrg6mPLAKTL5HY4r/uVrNjF4d4
dJAtThbK6xUdD/0+eXnFJMBDTk34YqiAmcOsRo49xokVrE3nff+/kMlVTqhSe+xSSFq93BqdI07R
7w9DRvxuAxDg/5MOSEN6Gk66uYuaj0itQnosyI6rLftD0u2qBp+N4wElvfeXRuOoEQKWuyAmfATS
hzqGjZ/Rd67RssWS3C/8Pgy0RGXWQmipeAlPV63sV9NewNDP3aDgF93W/BMHqNLe+Yt4AnoLdRG4
Co170sQGQ/jaRgjE93PEBe4/s8Jcjm2Bk9nWLLinIoatojzAmcn3F+GX9VmHRm0pXm1JegRDhiuO
zW5AA+Sn7YbitQRtXzURMMrVmrt6WbnHFu64yBmOHv34hUMQ1ZPuyixvmd8P6UA9FPCawwEea7Em
J3KQJIbSy5Bbi6BvmgW8o21sCp+ZF3x3lpUdIXcTOznELwNGST+PZhqpTV/fhpiJlP3GZkVitG3g
vRfxCmt47/6cq3NO46BafrictUt/sEszKnIyQHeR0YLWZaRFFvvLbtTadi/b+TlIcPQEE4Y1quSk
YuH7RVdaDVVLda2OljBZPNzEW76e8ah7/WY2+0/0PEJ37+blDjJgPwDhz1LXl9tSUSgprXx2b8rD
2z0/kxNKiFaVNAoRvSMSbPnu9X+pHnvLP5+2toBicho1LA0CgyZCbRaBetp6zO5oT0EjH52qG+WS
66tEj6vG713K5+DZ2/25T9cB6Bjs+yEWy3avZoknO+AFu0pv1lt/iSnGTJya8pKvXks86z43qm8g
NcScZtksA71mWclijpTFLXjcZYNyBmn59bvnASyTOH1FuC1TUSs3KNvc+X6ssXZH1DqzqE0lqBCg
3oxIv+KeYPdLa5vrcCS0TuN3c93ROhGxEiHRoyV1ecVQ9u2n1HNGUq4gBlzasiQgcXJQmbj9gnfF
vjIaHC9YKo6FWbifOqQyoE3uHDLS8MHMcKVnEzGyjJ9LnBKlyLbiGbBtBTr1SM5bV9zip9EPsXOD
ec2RvZhbtVuGZqy42HkwxOZcIQhIm1uxFV3t45WuTMcmbKJTDKSJXl3gESpdaMpyWmJpBOTni/uX
Ur8ayRBdHx2aLlrC0Q4PDWPoOTX26v3Iz/Ku5mVwaGcpCIlnRkUrMTVVy9x3oaNbEI87Uu4qDV9d
RufSUFmj0RMYTIhFEbZ2pa/480bZeTROuEF67U5cDX8Rw8r6+9IGfg/7y3EISIOZqkmMofHe19uL
OP/NMc9QtRfh2dt1JA0ioGFQBC1LmxBUuRZ/Ws6RD6C0cSrpLdPx18sDvq2U7AnhtEc6o5SQDHAE
Q6WlkGXzVEqt/frmkCySQOo5iHKD+ojZDXBDFEpb9Aou1cdYc/yHdI+lNJsEbAwCrrXm4LVYp9rn
ePaUjpxutgTq/YFo5YdN2Q8pO7sUEbmNOsUv4eR4BkkLtm8dBndwPx29O72YP14ZqiiEk93GZ9RE
I6Yyqo3/TpfaZQmZOxmOn6bTBOzjAPSUR8a9+7cO8iU+QDvIujRSN68f+TGc5auoN1kl4Ll3SbAg
afgNs3dIOH+DSIQVsfgmEh1G0h9w9JFuV1LxxGF0REagwm54DhgEQFK7alIgWyz7sUqLqUwROf3P
munJf3m0vdIoPiR1WNJEvnYtyswy/qBeo5G5azXFf4pEYwlJUMeVNSmNt5ooMcJ7E5jaa/KDHGDO
E9ykj3ljramZJGVe8t4STHnUgui8dlY8+upolk8/tKVUzjW6XuZy1DSMLAB/I/L/ekVKYFuH50sH
OVAuXVauugwv2XsC30JD1TMJZhBFRU1F6LsHG8+KVgVmVV3wJvl4Bdu5wEnqBaAgxCjjKhPA4SeY
CrwU+osva+MYG0hxelHr1uiP1DKX+OnBvjQqliQLf+keOdrt0Y7gbVqeIRCo3/LvSy93kL5So1oq
bEcGPL3VMYWq++RQHO5LIwLs7+ty1+bzDs5dLvnpFbHpFnXcCmeZEG+vH2UTDEzY1XFjyYP1CEb2
qJq+VWHN00bxs0vjg9+pWMRPJa1SPHR3mb31SVRwrzwp7npea3QAaNWc6CyZhnzSkR0wrfb7JlYu
nHvfEHget89ej5hP+bskGp+7hoW9V+jp247TXF106Ayzhc7kGS3Ujet9/V70hGfFoyb8l6VKNxvL
wbyOe1xKu6OTw0si9ljSpuYhMVPeVrlHzvii52Yv0ml785jz/2XkYwpJy4T5hgvnhMox8Ed/drfE
cQG3dHVUNHBnsw1aq/VCuIbQJ60763uWzZYMFDB75Norlf4wJigxKsvh+D3H2z02A2k5bJjAkK0h
QpnjGNqcFl/X0/uNzIi4IdR1oDmV5EZoDA3596Z09bcGDYY53+u+mKKHDpsUYeogGtrWvuqFw6s2
gN9NRvLES2Ip0BvYDhkR3+/m1YhkWnb1QVlN3hCynJ7rpMmpVPO/oiTv09vDvnmbBuRXyihtYlch
2sInwZvyfPiZsjnR/X1dVKX+bi0hK07RfRQ30MJJSHOeXr6DleQZUKm3txcnpZCGUHWzrIBUbC35
7TsPxH1QYAb1qA50IdFIb6XhiBdZF4Jw0qoytgApR6r7soaBQyXBuv8Bs3//9W7VLqS1mUcvr5Db
9tHOuYfjEvynr2lRm6+HSUeq+oha3Q5sZkdKfUtnzSxqSKtlJNEkltz4RCbjoIE6UEZechDctZLH
vcNr8a6JSxwgjnx8B4WmhBHMCLfZ5ioWlB5rH/XJxGURitDsmSr/g5/UYmev8ltMAuwmkPeFu/if
iwiGyTDI+xL55dRYZRrMEWp9dDUsMXVxT247sTTa6KZxfrKRrx+PSA7tisA1pL6vBeG5P8w5kIiW
9QzhTl5OcAMaFfyb2uBOMU2x8LtdPirivtATLqDJMlb0zFQAcqsrE5/HBYzb/aUJtDo4sMrf4H18
KiaFbEX4lFRhVD9ToZbWAv5DPQhDQGb9yxjkMz8moEXqhT/OnnLMyqOCtE1WldUGWrCJO1t1MBe1
fuzdCw9l+RxiyHF33in21Uj44vk4ruqohexoJqRcYYDxneLTSG+v0R77TkYvgrSpOAPdKXbK/Zcs
ct6TLH22TSxXKybez0Y2nZvurRQKtqCN64o2y5rwEAllhz17AfL5wtFoKeRUoz5rPRKVQpxA/Qrb
Gukq9UbywFUTttFlGZjOWulONWsIfmNdzCJDz7wx+/I+aiHjD3XrUmhwv0X+t6gDkWL816kQGLnT
bMZqaqP5o/ptFeIVcqL3Dm6nHTUyu44E3P7BMWrjsCa06RlSQjHZTjjvRwq7Av70req4IToqUvWq
rmahbVMXhVLEAB4dWw31VaMAj/bhuoqCqyQVaGBXN3OCMlQTY5iAUMfarQT1FePfpy0sQZ60czIT
pveOEAIvsushI45kY0eYhVw5TbCnyng5geyBEN0Tzx1GtFw4wasSbXgnVZNxXKydkcT8Vlg8Hn/t
QPSfxEYIT/iVyLcsFkAQ3bnIMQVfg8tNObQXaH7dsiszLVKWKyfHPyLrUifhIqgqOCGKX+XYPgPj
rn3R67ZLFWg9fsdjiXYqYlixrh5+I3X2viecwNiVklfQUphiD5qk55LGyq/0RdYXuD5l6Sno0+wO
5PAP7jsdcjubgwEtkg70mHquLwj3iWsjC1PMAN/NCuMPnQeQvFDdz0fhRTp5uiQkorW7IUd5PaQ/
ELu6MvjMwt0aSdXWOV+H/uPB7UZJltgLft/dKTc3jskRr1W4OW6iqIcM2YhcuDQYKxVLq5+pGtPS
qO0Jn7bFwNpUi669wxGMaBcy9Nk6yWNNX9qqEix5qxzqY6W9MT1ewHzcRvdCuaJx2mVc3aZDbkVE
n/cRHsliripAFivKXu/NMllF1YqOcqNaR0rmlyGdQlCL7Ee+T4y/Z0fkuuT8OcGcU8LsvW9haoAS
WTjxMeiB2UWKOOKuC9Y+M+yMSbTRBh7Bgv4sZ04x89vM0YlZFP/J6hk/45vIsv7GbBDs5t4iWotP
rPkLvcFdlO2F2sp8kJozT9FGdY9ZKBI+dRsOBBffO9kJLhdWB+KyFU7DBQhc7Pi/UtNuvEImOK72
kZfJrJbdJGYzwGoGmGzXXpJqfGVH57937RD1hQuaAaAKI/4rosGIVDlqwwnBcdhFXoXW1mXFFy+E
lOKwDQDit/4WGER4hPEWjJo+khYH7j0I6Y+WavQ7CxLKUq2od5cZDxcqg0qfGgsu6KOW6ox4d5ge
pfuPHmhsFCqB1G5qxkd2D11YNHH8vqMl2cgxL4X4+NbJfmMHhyVsov5cdyNo5iXl2JupGxDoFmAU
p8+FjzdBqMofP761X/QKJEoq7uEs5vdV6OStHhrZENaBFaqnj5EO6Nf8QBFd86vMuuIsuzTyZEnJ
WV8KHr+xl5d9m1jhlmiHjMs8FCGOCz9l45JGVh0Q4Hwd18v3UKKPW+e2BjAMhYbXVENo5OecRFJs
O9yGtga+vm7foGBDqrLZpFYUVy6gBCXFt8Ps3zZj8VaB1GwZLwoB28pJGYMIga1yHIS9A7HklMTw
6dZ/nnf9eAAsOCILkXadon2jIK6Xyo33WlQa9VuVkmGTAH/etiCgTpO+3P3pBNkc7O5yzU8vAhOm
Zl/uXrP4pvlzd7CSBPAOnVoeK7jNlClI6xfTXAK0JohNxLgSmFVAUC7I6k3fJzZkUmZ+kPNxAYkD
HmeA1QWZMx7sTfeU5er8bkZX8l+5ub+E4rbtmcEJ/MiRb58UrQYuikkfGvM3CWLGs8S9lgzx+13w
BkF/xuXGE6VgC/JBe55GPFTGry4x+Bk40eCNOsZ713ifjPrHLk9K/1UTEmIGse7rcsW2SvFE7s8Z
U2BE5Md3jS1obpqkwu77gpVlPvP3l2qyuDl1kTRXNbLCR4C5SRPSGm0WwncDWAv/VFQiBMlwCxn3
U98r8QNcWi2fY+6pfnHjnbM9aoQvyD6Wz+0YhmIEwavGSddyca6grBNwV2f5kNHkZcOPOGH//0x0
aVbdeU3QABys3NQSc/xOJJ+0WsosF658lMfT417MdrLxYVq/oV25tqdjM0iaPYHXRv/Uw/Av4YFO
qw4JrXiiGy4THAmNcfQhKuL972VVgUTyWFUjDQAi8sNpV/JCJCv5Y9JIZjL/WvIWUxKLHY+UDhod
4KWxgiTNmu6aAbgRkO4jWa6bTeGbRkYwn/rlShACTZMGq5J12x0psRKBiq+me0ahLENCKcCqXG2d
xOt26G54rZeQ0Q5KfN2sc2qXGMb0A6K92zrknvAQj8FhrJP2xFeWpV4L07LKyf7XaejenZKT4eQv
azxsJbtAAvty+vLRH9cSEfTBNvxVGdG+1hapRM9iXJ1GEvaamTBWZXiACChp0aAEKpZoH9TWoSbk
QjnrDiWFItPVpAfFe3WU9qUu0AH7jcI14+7UoAgMpmqzUUaXljLlSIU2cmxXyLojxJKar/VIghgk
i8aBPl9u35jsXvQhKvzaTgpWPZ2npyaZYoHpWDSLqr927t9XBkQg/KK5h8UYE8qFTgnbTxtkIExv
dkZA95/IYtgVpL59qdqHJPO3/3hSrTo91WyzFMrYlOB9Nw6pklhs08E7NzNFR2TZ4EvGX7HBfQ/f
wnPdrEVMcJ29RC/ek9owyKAegzwk1mlb1PdzBhhxDrj4e95wenkpGbbN/kqQarU4q42ze0QI03Up
x6y71sgNngWfYTZ/yETPJy/fcztDsphQiiT6CLHuEZ28esvpOkyRcjs1qn2gXEqiDSqe9qoxU0r+
iLziirniBE6MyV96yWsuUCRmfeCNAV1qKaTxISXWU9hdBgYcK/MFhO0jGvp43TWs+Us6IJfRryv8
zM/ztPxUAICO7rFcyyvkKMIV7y48PeGNb4hjpWHesRCdnuBBkXJ0O4OVbGKCXb4MobilEsmSu/0a
DAA5GEpS1ASxmwZToeGargkAbuRBPBMPzOJmkcj0HtgH91ZEEdevlCtu2VR7/IHwnoU/yuqaK8DW
24WnELf8seaHxcodBYn7+C3dFvFknPGqcHKw6ASBIJjer90LPAVx+uhfGST9XlicMeM5fkR/KDKL
FwfMjjDdR0eC8WMoboH5B5chraRjJOYIul9L+Sj1u1dYP3Dj0Kjwwxbkvwxx8yEezhyQb63yscOM
4UrZtznX5Kl8JghEhGg9zPLdaOTO0KpQj5yfmTZkZVLIqEN9f6DlGxE+hSTz+dzW1COqedC2VVkR
Ozl23u/OZyPdr3dUObNDlgwGVVsjZqkXdpHiFfc/js7LpQ21VNU7nU17MYb1zdytt8GwbvRurzQp
sFxITrINK7zknNrIEgB6RepP3M+ZQKOpurPH/NI3wQ3o+75ATR8mIVfX7/1nc8KtALsck09aicS6
WAwJnocNdmDEdZ1rTDdGv0jJwGg5iSandilgKopIXK0VyVTl+yT6IQiTeaGGCWtqbTjeFwxC14Pn
NdVEHHoCfFhOKgZulubozsxg2RhK+7mvfqq4mRZDBmnB/mU17NKS/ozf0XmxC/nZ/FapWSZL0MzY
7mY0DOh6qiQdaHetdrk4zNhkPqG/3hwMzDtnonut0bU2QR0JPAV/HY6hRm+IgO8vkdU8HrK1FBjC
EH+Y9UAzimEK3LKNSfu5w1+zLTdIuf2XshA+k/TIWcPMpizbTWwAjop5KJDUPFQZjnTuCFRyRgXJ
b3uQ9mbuVBRF8CYquw5+S/tK50l8IfY4jvN/29fyTGg6aYbT5wPyF0uWdG/NlKBbWhuX2At9GSCi
sFVqOafJOC5G2thNZojcquIsnMycQW7XjSEJILncQZgI84XF+pOu2UHhzbxEYHXRowySk9owligd
yOzuE5t7kMYTKQRnWLoTc6CIA+HVMn274O+RcU1yHlyXjmOut6JjaydFNqGHFfdtti0AM06YyAFn
4YU51ikPGBs8U9z7+EIVUhU9m4CIVIi988mCrm+Nn3F8zA21t6oOxJ/9f/MGX14tcsLbFCkl62Jq
ABjvKnlzqm1x7GKOcynDBa/KZirdGKKV9rlJGidOalE7q2+w7OzEFxdwJCylNohhQYHYsXAu6P94
ZXf0d1UiSVQKfGfV9qw6AMF5tgMFs/HLKmTwpsmBOca0koLxCikXGznPsnQM3RJiFCwbTGVNEnsO
G/NYyniZZWfy8sWVGEhNIeujlcN8aCDf/z2qkO3KCSOUtwhY9JhoyCWyeYghlhyFFLsx8bHTRQ3k
JG3c36/7Qa83kBIJsLT6c3n/x+gnD4BCQUfh2AjAqDL7DWXc/P/8uPhpiebsLBw9h8TskPbqhzB5
34J3aTIj6BeVx8FqUIoC110irWmUuONwkNQx+VQG24XbXm1D+Zk+Ll5shZJV/pgGPs4c3IqTsA+V
R4i9QAu4SD2/QDZ5j52Kvvsxu3HMOnNE4RWpn/69t+HoLxb/x+mtqPD6cfOyvJsBUYlYjrtXJoGP
Fe+/J4zycqQWmWSOwCn8CBgmC8mzPTCM1dUXnDDCad37hgPe4ak4zfuNTo669TgktnvLI5jArHSR
WQaN7p3vF4m6jrR/xIPHQLckjJONXtxVqmcqMeyxxRRnJsFsmLAG4eToLsFuHna0GJsVD31H0r/3
ysXa3GREr028/AXe+L9sm+euZlsTKhZ6bTTuSPJdxgTHoSrvHRwtoDz9QcwlLlBL7ls26AWIkmuw
hayooFmVf5iBci1RB3k25mx2l8e3J/cZqAncplJeueH+UOFNtUiY8SYylcUlc8WvRRdFeusfOmeR
yWG7/qFFtI8MDVsR30+yGwIgzpyj1zLZYB4cg4j5VhA9FtlSFYn6S8xd/rzap3rGPF1Fq0zmVf1g
yb3Tkr9EIKCZyATfRrBwX9EUB0dZe852/1LqY1FZltEXcBWcuHFdUmUd3ECb/W7jBmtRCNgl4coc
k3jYPS9d4DmfA/Kx0FruvAjKoqHqjH9Xr1JFeHaT16Q64CxKTDAHe9qhqqgkPjC8TWoTZ+NQf5+M
dWDi1uYMaZqQXvqN/rKaaQENeVvFfSTH773gfwB3pOrWF7AR9030Gl5CnfIzWYVXKJlfqzeQdkKR
KBIBdRzOoPYLpWVoHcsUL2o2WiqyQrnb+uc7UFYSoFBdZk1AtV8Ji3r0/2zMrKLMnvvMDhwMrahu
sFcr6a85st800Cv9ZzkY4w0o3Vt4Xw68a/2aTBGD1CIbMysM+LQvwJq9Gz4LgFv570QnVH/mK9px
ZrCYsf2AqbE6WpEl7tb1ejo/+nX0ug8KwfNKN++R56E5SXgIHm+KKsKiGxXoPmIu2zyoz8wqqfNO
f1mxvfSa1ZPpfQOJgN+E3zhpuDkxhQkWlTjrPCtpjk1YGU3ACRptaAIaiLI+O+o38rnz+DvvHJzg
WV049TWuiNaguf88Jm8NkK6hbMN5Bro8etGkWRTIEfi/0xJgad7RB+YnIo3mGCRRqxaKXg9eK94o
x8qDSffvaQ6HeXgjOltu7nlSooGNXrryEzsUQ8rL8Pxi4npSwE0ONkYt44zfIQAWT7UIzbAh+FAZ
LeEE0NRxUfHDPHMRlOJOtggKx53lgMQoCuKYWLXPZWPRicKd5SATLEurZ3hu7Bs9RRsa31q4ufIw
uy4OGcnk8p6KOJWGTLtUhFjArUl6lRpwrsbfIB6tycvmrngyr7eqt25lAqMT7XrXKB0cOosxtIIH
GWdSSdaGbH7mB0XjPDLo3/AakFhDT9me76asPx9zHxZV65sYLZr82jZJyP9RfTkEOeMp+4yGVVT2
4wwIRGB/+KV3qG2Y204/aLPMu+azJFRDAkb0+O5KyWEFOPT9yQG9TV3sO15NxYOcuFd4682zYIun
QCgdfNPpj+q9zmgmimh0y834P3mO9xZh6LllvEpm1fIsW34dpolh6A4uvnZD0LoSGlr+6PgRXOz3
bUi94XtuIKqnQt8KA1BIlSgFUsSLbZvvYhop3uEfMyeuWtzfcbwqWbHc7oLm2qZZZT21hxlCscml
PeP2er8tdM+hus/rt+bHKhdTml7hY1yvK8d1nXCnbH6lo6t/ACKoKkv2XkN0cnhXoBqttQEcNMSn
TcN79FhH5mwONMC46KvCIHUIQcO8KZhGzTDlS7GuIbg2lXT1EWUJ5/T+tUczSwUgu1gn0UkJffic
t4jAo1e5mv0A0gxFm/apXhWqaLEyS/g//Xbg0lkDrEUqSi4d7zVVusByyDuOSUmL79mQ6Nncktii
qnH3WaCSce+uPYM7Rp3gAh52DXr27E/x756oI0hMbSBgIsbSOTrzNmbVX0eGbjFvJUvrDBtaa4/U
HtLZBPN0vDm0iwfYdytXlFNA6ZZcbiiPmT2/9I4PNbc4QVV9PUqZ4QdUqru2RXxsfcAxo6w3eu/t
+H0S4qbD5ov6sfN+tMvvjzqYsNvbdJ/m57f7zBD2Nib2Vw3O+V7W40JroEpgCHZP9ZdVnebpirW3
UWY0yL1cW1G/neuJpaKJYIc49tkckYMq0U9SIEQhUH0sw47wH+foKOC/VppFF5ifLUSPYZSLm7TL
WntRqdzb2F+nBxmypKr7IKNG4/SQpAGFDex465MPF6Qn07ee9VqpNJYA9HObHKvNgcgMUlCgL6+J
M72tbxRSkKDJIEgW58QD/NzyWwG+mNui0XFma/7pCvkcpNQKoUbWzUqLnzVHrGAXaRLCr8kYwQGz
Jyzm75KsemyE5Hk7myElfmNeeo1HxXM9fJGa9Hed5hpv2uWkhFI/kqJIY1RKyaKx5Kda1gaAaR05
jRSYqWxUbYMWzBHJaA+mZpzcqiEcywMoEHMCu3nX0x7p7talzqQmGtNai1EmarsKmOxFAivCncDs
c7kFqrlgZzXzalLX2g3oh4XDrTKDg7s2EhWffqnLii5lONrwEov4CeSML6yUT45Ay21PE+te4IeM
ZtjnLu4b0t5G2iMGpt63tXG+r9MZmNzBy03DEK32h7N4eUkY7SjqlMCsB1nTw/qsCwD6vOeRCG0G
o6OBJYUF3PjPEU188pl2qdHrNrztWuNkBA43QMXu6YeSnciCO9CatQOctzhYU97/9YktTFgbuflu
gQbnDM04g1BqQmwfir/b9SxWhrTFM2IetxgQ4bReQuVEIg0KTn72dfitn2nlP0eA9wB+hsblv2yI
KbjTZX2qPQ6vV6j591kCyamiBtd5PB4KnSS6eG5GiEqbzaK4ZilluBJfKEXK6ClyEv2GkDcxdRW+
t7ZK+NrG3Oix41rHOqDXrWxrXKeAAO+4iiomwBSt5fP4jImX7e4Usci+NtDKRwPSnrsrvHUcJ2qQ
UOpDTsq+YGA9BqPopYkfZJ2xd/31po/pVlTHDVrgAd6WJKfEiXcCjbbYa/ACwVejDqEU8i8O+/KM
BNHoEr8gPCOSrU7G36RjzPlOSFVgIlg+ANKOUZjJARSjG0CWF9hX1zNMNb1rcLUh4IgktUBZdE2D
g3cbxNimp5914uQVQM3CKE4gbGAG6EH2xrwd65zt+oax+EyaYzQTDYi4KvrOtH6CzYhC4KSWE3OZ
Oz3tecwoUbD/XKnALJxDfbu6ZyYnHZeFGx8hHE8rQdxYMJ97CS8dUn2JSYWFG2Y0XGX9CLdyknhP
SGyv6yN2G1lQAuZ21CXBDasLGeFZxHSKY3OiT22OuKhxg7OHi0vl5J0BX5BOXAiSlArBX2kPMtne
a6Q4CRaoaMC223JQ760VJs7x+iakucr44xA+ZqwztSXx7tiwDOSqzJE0ukm5b0Fb7MViwDd3O2v4
cL9X64CwhTYkqJJJKRegAI7YSmnGe3vStzBSAVjtTjnW95rsY4qknJQzOXFa+DDqxlNgF39MWD9k
jeyVtZ1b4XnLGNnaFhS+u0LTE6i7ZnQkFY+mIgXJVziFBA1av5PD9+GXRbij503jwgzgABStVQfz
1nuF/ZBWGcBIdJw/nuDxJbxYzlYN/MAPwj75abBaM7z+BLxylqJjveaa9NR3OmZFrvLtLAWeGM7/
V9ggwWS1Mkluqf6FDNUn46zFKuDVhUclwnZBz4IdftDXlIsrQtmI0FL+9vsF7BzY798hCHyYDEqI
PrNB5RvHjtMICdQzUnFnSdkj0Vim00daFRF8ar50TwlSccxiQ6OrH21CwyjVfAWZpgxXpzqALlRl
71y58ZTog7SVm2NJphCyPFSvKq1xCUG28C1GHkxd+CvYxrSd/NjYOTDxiS7pFHCMnSO2vAxG6f7o
eIH4kEtBu6iTj0QQE3jwVbmI3qexfelJ8VtcAo5R69N884yy5qYJBXDxV927Ad3V4IrynzThD5Bq
CzM+NwTTtu/SllYnuVRWMapFsaQ/UcJlTtukA0haAm9Ghg+BRbL9mMDtV4Wjk5mEsnxfKtmAkVuQ
uHm3ebj3u4CmCEIgveUkmFXYPJW+6nCFiAbhWCBPnxu8Jrk+4E+KcF/+00nBDeFRamPw6y62EJkN
b+FvKUR2d196JN49JW48CbngzEqXdn15j2AWyPiTd5I1zlQ30J/uK7NVOZBlqZNHf92ygEZ35jeB
DkgELMBCX3J3b2/TWuPxYgbRm4UZS5ObJS7yVoCqdSEh7Xa3yXOaDlo1VVnBODrB+Wc0+eO9BO0g
SiKIxkFvBvE5jQNLYIziADapNlxm+Blt0qB8ZcCmnsVjlLYIsYQmxPYqDTXX4avkdg9fVgyL8zeF
DfKCqDP9bZKLwv6hoMgs9W/yqiLIQACVx4JgJY6GnG1cXg5XWybbeOD94yuwOFk/5cRbQzoDp1rV
KHyYC1DtOsK56kwOrVOVlLvj9hPuTWqXaSm9uNNxTZtRXg49NDJnmPyKDjcpFqPaumd+o0XBCBEJ
PKnNlr1oT6PoxcEysUkw6MtdxujvAZYtJE3fFPB44+AdzhwBN3A14Yu5GR4dyDvk0w3zwzkCTFaQ
J68LR6CwdiI3PhYfuocMm0HfW807kV5cb9YbNd4L5ENfAY1rUQjE4JI2OM5/BJwAp6ROx2kWiNfA
ohwTT+gqbPdBYMMXdPUe9kHglVyRImZUFLhDZCpiSOmebLBCwj+oozrWH66p3EMBv7KVxUg7VsMU
HJ6wfo7hvAS09lBssTTNoxmnoZuzGpJSWclvPGhKc6XippaVpn4nY4j2ywN0WowGWSjKNAcVTaxZ
SCDzhbzbh+z+mvq5C1xHrQ5CHayWJDgNR4yJTW+jTJM8+yG3uu6Dd/89RflDBcQoBCY5OHF4cwwV
P77SAwcfenfjCGXGzy5nv8ns+ydUkkdnpIrhbBA5Fhas76odSycbUPZYX6/Zt/M4fbTJrVYz4KgV
Njhxx8bB7bclzzx1lgxYO2fxhafjDL2Z/dJ76/PtY8Vkd3HTrW8VcrvS5BvZysEyIDmnVEUnoWdq
o2XPMkM5d37Z4YD/oit9FIZ32cGaIcmXGbsqoOyB8Al5o//WHvv4cJpUmA9KR2+R3U9XXlce95sV
BYzH8JmtMbP0TJhM6xJo2tq4fOrBfIPbILsdpXEMQhTxQBkPsLmJ5LOr6RFvBNcU3t+H9P5L4JMS
CLvFvLriS2Vme7BeeQrOIetXmFFOicS/gfiTnBfjGZqohagnJhaNhISJS2dyNEpQ3fQNXaXa2/UM
sgnp3YOSRfNtB9k63pte/OvESNMKqbQuO2FNgQN9fp9Inv/a3dfogcWZRPzu50w5xvrq8sd9VA5p
u48nGXYYhBZqgAF27qH99bobsd2P306tle782hJC9Ecmegme5sM/hTX0oTKyPu/prSezqXa7m3vI
m0LQxkrIU8tW6FQ4a0CWZgVevvpDPxH5NKae2PnT4EU2Q3lNI3zaQCc/YIySfULjI3Y9hfc+ln7G
gCgLLOFH+JoKveRcpMfXkLhie9Cz0g6snrU09fERIBlW31XfXkTt2VJqJN0cT5xdSHZ62ncXbzFw
9HrvB+f+FffUsPxdyp2axFP780xCydq7p7dsGIbtS7lc3gJwyS1Efsg7jL9JoxKUBkluXNXsukH6
Ci9RWDlQ61dQSfTqCj/RYm+28xJEsWTHLOSy8Pmk3nd9WVfkhaOT6HqCB/Q7VbCS0FuRQvyZFy9e
xecUacEmvKHCX5956ZrWizXGL38V0lM7swEHHB+QAlfBmeuGD3WEArdg/NdEMD1gfhq2M9a7x7jB
FZqWgAsPy8JnpwyamR1B+i5n/C9KwtYE03ttkozz/awnLl53AgC7zkinnn5V7cJM7YR0ZI2hOmBM
xLvsNsd/J6X1gqIy0sQN201xk8HoGWDc88fFs0TYg0617hB+ibdhRKoV6GQBzjQjNeX368krZ8nG
dhXxNkmvQsTsweWVIWwxO3TkFAhJYSw6TZe+sBYFiGFLI0yd03kjwJN1IMFMxn/QpDVQDKQTQ1z5
YjxUCL4XBWFznQI2xW2bJVKlusDzWWW8vQOqc03owpcfHFIBCJlOh9B5WqSngEPhVn67h5blz29c
Xj1yeDx/2gS0HnIqXNVkd6rbtcOjd6vvGUo0TH1n19SSd6Y6c0+nNZL8BquqLyFR+81pCgOhCV0w
z3CcNIhUqt4cpF/5DzaONAcUF3hz263Lz7H5s3j92UqMHnmgfIbwcbXGT8fafvn3ORfUH/UJt6wE
+H8RiFXS3oNVJXU/et3fFxGm9d6DdrmKSMKuWXZ+Pns4ox3Nb/eGwzJoGVwFJREY8AR16OBySr/9
1auOtWtBi2lbzN6tjGWE7Gy0RIOTOAJ9IK5vED0C7M7LJ5AmsdrJddu+HINyCfjWDf5Q+YMCC+lf
y9PMyIuqRVW3WOMnHJOuhW4g/1HB3xwIUH2mM/+9NjAFK+atsHJzNPFhK9mJJUiDlw54hy5ERxnk
8pKm7fyMru75widadf49bqkU1vRY2x3ylAkBGhSVzTTmn+UYKXqj1IlFvPuw40xYfDeglylYSkFy
PtOoyfD1nrpN3v2BwLx3/pdq21XM8AOfHS+s1hRrFNr65IAHL6iV8gBwUK1elUhk89xeVobQzgvc
jvVlOUaRe+c6fgTbv5QP4EyMCFX3BLOBLZJf2W7keKtSA6hR3+7+Sh7tMexMb0DdzmL2mV05W1gj
F73NUl9Qv453GVSepHmWGZDnG9+G36m1HbNO/hueOWNdL1iFuTqQfs8FA5TJouaExxIkSmK+06LC
N1VEk9CRluys2FCc4GRgyFcTQHYtfLhctmAMaHC2WJE4Cl8bTr1HATNwZWh6xQjM6SOQJLbAaQRg
pXfkc3cmSlQySP4QU3QQhy4LuzWPJeoWZKLpdT1ttT11v3kv/JsI1a5xNOIh6HjXE49OGjZFtxRE
kOCsL6eqUAIUgJT1KJI91xCHNpd4caq5kTZn+C0FEwCv8YV2TnbEq//LOMB72WWbwxTF6fFX23OY
A2jzN/1IB/jixYzmPFSbVqdThJAEakkEH7mFJ/gy7ejO7byuueUNCMacyrV0u5xXZ3f82SIyVaqn
DIPArRAH+nV9QqzLGP+05OqCaj1KSM2RLOAWPUBPAZB0sqLMgmiHuZ5jwa6iITr/SHOvsb9uldVB
Y94pMvIy+tubOaPNH02y/pVGCof5LUuBmSOd31+ur20qDgcYM8OrYajpikporDdF9ezLUQPPbzFO
MkQIQeYFQ1fa258egIbgcBYjfjiWMCLi1+OKt6WlpYIK+omN2wj6vW7GryRLTVLHH1GQZ76naSbC
Ygl0LRiPSoQnbHEPynmmp0C6bBOwBGD8eKU523LWT4FovH8ClXfAZVVey4UhmwZDjqBXuDcNUrAv
9KBP6Ggg/qAuShcs1B9cnKZWCf8iZAYJCo0FkLKaJd+FD4h0ikqQj2kGHSwAWOYk4jUd5t4cnY7W
3mizTGtcx/AQ/Iujl+v+cArTt/5ik2m2D+yu2x4GpmgZk05V18bI71JtJ2wQxnqBIMEtUahJaEYm
rGSd5HEFgAh2nSAUgme6GR0zJ1r0J3ppHZVMnJo1EXX3ck7Fe/CJBu45KuvvAFEElOc04nmmq51C
j4xZqoXJZDN9XSi1hIFF5V4LhjLIRT+xZj0EpKHm79gCLKI2lhva/ArEKNF20oqAOi5QsKghiLtq
iEOk6acr4dj8CXxZ6U6ET4TaCRjy3zxHyW6I+XJKC2dcPCjfsd7mv3EQauvtmM6Xx+y7ezAaS3Lf
Czw/B/ergQ/kjrs3C3EoS/hB4lhYahDtpEnxcLNuXneeccNNJH2T/7sd8n3+Qd7tNmRNtrhWUCh5
qGFN1PHfpbh6DES1kNe/71emjzyQnHMag34IJ1FeVeuI4nCex6ichYV5oGTLKgzlXoLarFYwa+F9
4QsRLd+/whDhglMPz9gfiGxn9AieHTe3lEvDSciV+4slMTuF7ol2e5B9djhTluyDVD4rTwepkBuP
mhFqcunhP9T4p+6kKn0sE43gduDHJ8WuRZgAC8cxaQOmugZzKay3k5Efhg/Q0MZEcBtUpLwJ1MFb
2ttuL90HxV2aJLso73D1Tur1MNcQPxddwaqNQltA+sLDCXiifQpBQE5vtu0kec7x20xRIkb7L9ty
eQZTzZZ3ifR7jb3TWyeOqdJ3ggloHJv/N5oiCAmMpm5xtxZhn2JBmpHwrEQ0wwSJSKtY+NyWYLsN
y0/SmNjGhLq8biPH79yvcOer9otekoR+iDyfOpTstePuqE7NqP6Z8/Hhu6x1iBAvz4VpkZ+7cyIw
fzw2DaFhzKxe+3niSKTes9u9kWN+Nw/Q+EjjAo6C7jxXPtp7piPNp65WFBH5qtOhYyLZ/mEFStTe
IH9KBnxkWT8DLZHCMpG2MDiLQWQqrboNDgkIRxX+iU5hCxkmzL5MvvlwdQgahCsZXWhq1qblJM2W
wPWfiAyqwojRa7TDMTlRh4RCLC2vU0wQooDSrzwDz4NnVTTwslze0NGie6Z+vlWxEblD1sA9DQkj
J2B78XE9LYLcYIsLDcsdklD2HVs6Qm3BneK40cfOBkMnHidy9UKsH4qRbdEd49C8tDSM6zrDMUcm
aeCeMSM+pMdLvxcwCmFmqCxCFCsUng3iMnUFETpF7DTto7pWh0LkzK5zHIewCyguI27wHeXWDDA1
RQ1IRamU7uqiW9tFQ2orHK98h8V8KR4lKGK6lU/KJz371/MFHFeDNXzyR+sAyiKHPDg7G1MW9LGM
ovepsJ+OBMh5rCTQeaVyfS5BtvVuz0+NktuyBRUMeIAgfSi88lHYN7mVHgQUGEFgvhyqychb8Ys4
2OzWBxhczCxTYFU9sYQ8u2wKfvs28hGc/0/EzHGHjwqnZo+qmQlGJXBvGRgaRCfdficQp30luMmU
iEUjW1V6PLxY1PtdHb1FTFds35SEHWiWaTmfSv9y0BHdo4j6OQ3ogVzejUJyeERRwOQywo+V/vba
WBGSHMlfVNaG8MEF8e/120MNnIAf1IAFr4qq+4/SFFq21mzRA/rx2d0n6x5l/1yoUGcn8nSZXE7S
UJPt+3CbGJbdjF9PJdhiqHI57hAnCL4oOV+7sBsczDG5IuT+i0bY21VSVgEkZy1hfaBg/SjQ36eI
xdnTXULOKvypx3UQsnH711gOIU9NkTYMkkphFV6ePOuqbGKS2kYIybzud9+U+HwSWkUCv6KECu+H
md/NIG133PyTg7N+1c5UZeZrBEJ6b6/DN+GCWoB1qoPvwo/gVxdKk8JgFX4+8gBbTgLy9Oe9jq9s
mqfn4QbW6er8R2T2Qyfx+ZMiGS4ZSf9L+qS5EpxeeUMKJdjNGoFiCOWa5UhcHFGfV1XegSYj9Ehq
jf96btNHhjm8VGET5jmFRbgdSvyyef/W3ratz0Cr30faGSq8BFnF4bPmjm8UZtG8cEWlrfq1uNnJ
3T/rfi1+oFOBw9EUqx9iWy1WbdaTw7NQvk9pIZqTsQNHfDw98TiKkTyCX/DUU8KIBBXuJpGW/u6K
1cOlEbhcwnTHIzQXG5/E2ib5aqxIhkGX0eyTZwYNMqllHULarzfEspIiCS02bkoVpQjom8mHqoCu
vhEp0bHdFqC7VkfdZ6yCcj7J6CwGzRA8136xG9amqBFbmbUxJyBmOM/A69hStvHEQrSAJ8XIKMXr
/HrdI60crK1BYllPkNz6tHEX1NA3qKQF0jfpd8ihTmHG73vhZVP/SIzrCuIsyMvQ2k05h+jV3qlW
6aXqLY62svd4oovNcATqeP13obJ4Z+kRfq2oPx2Pw75vr2zxyGlN3/mMkvibU7JaNhC/rihP1p1a
NZfeAh68UM3RfjsXr9n4zspDiAIC4aLbkIJ0cemFCvzwGNjM+6PAtcFh1O7cojsDyll5+eFK2Gqu
h6VLnVNrAAUelDZMfr1Tmjct82T+y0Mw4nj6IwlenjVar/EKQkA0cTvQxXF5btP/PVko9bMNUBeg
ZqjO7rK65Hx5295CG2LpfV+XT2cil6iqCK2c5U+Ehpc2PQfDRYMtdfCRvMRJnRjZbuuo7bzPen65
Z8dk3E/OAh6JrSUZQ4ccKLEKb6ZR0wq9Grn32Q5DiAzRuUkmRk7lRHXTG1RUmJVcFblnx7T+XWqL
MabxjEvu+1+Hq7fMEVzRC6L/hHUpItG9w0U4LuI2/Wx/vJr2j3kumTE64x8emdjqA6BYoj4y4shZ
kueoYHr5+ZuJ2sPEm113G2otcPJZfnI0MaoY07dwbdJ79DRWj+GYi/voT+PnH5b9p9KuK1iVIBZL
EGu6ziI6E9VbH9ycGWWy33bQ9kqHQ9grgXC7niBBYGhgtIJCriQr4lJOcpa7/p1tp9UDrkVvdFGP
K5k5DDQKUlI+4k9sHlBHuYSNsfuNf8YBBkT55baY1HUGVOr5CMJt3p8xicdUHezOLQEgQq7Eug2f
8rIA2EhFiJ01SzU4KJWUkM3h6WY83oSmUMSLC6o/EoR97f3PkTqhayriX3pO8Iwq4einjUt/qy2B
T4RIQHP7OUUHGAvjDOAyfkTBY6PlANB34YA/jIRzVUBBHT0Z4We3Le34roM33eCwdmsF+oao+iIw
D8HVB6mIL5Z3aVIoxtPmt+EkEgYt9ARVEx4ZbB6fTPKfCGUHVP5RsViZL48+80cB108zFldf6ofm
1u+PZwZHWK0FWYtgQ5eYF/KGecvbBGtPljPr4NuxvxoiTCumrFrNUB/rzW3bHoSEarmtu/vi0bQs
iTUwxTmmvSY5RX6v/kKZzJm4ZOv8zi79G20i3GGcukR8LpYmw3LM8XsNimnV78krKXUGVI2zxGPM
QGfiIRA+CEALCAFR/eHGvbg0XmCO4roYvraeLdCI2Ls02LVrHFAvCNuBZv6oYocshniXjzjbT/pM
+wcOyH1k39WXRkIH0EACK73jvy4rlYt8KzJ77mGMdj56G4BQWGPh5wOFNTNCOHLNoAf616AJ0hxT
BSGdlaF8j5YGijYe1GEnlz19ufDGIiPGjW3igjk2tcPMxE7QyuE7U3xVhFtP92i9meSKUQOf7kHi
TUzL7VuXkfwRgnnyvnR48k4b/UYGekTObf5yUW4Q76dG5iUhFxP/V/+xzYmsaIjptpPsVVRDOsfI
CjOybiqDxix672NIxYpo3qNHfl2XBoTtMoTFTwSp/utUj+rzL4OgE2WH+RYaiWi2sy0kAkl5hz2k
3uzzDfAHeTEOc/FpVcweAaOxjIC+2UBj1t4k6VpgOfaIher/6NAYuOpql//XkmMBxN9L3n+xI8dY
4qe4NtvwPf4deMOsQobIelfKGVwGuFWkXyFrCHVgUYKVdD5nsOu4MYZr5tDF6lvGLu5Xnga9Ayu0
wN4JjOlJefdjkswgCtPPFpG+lbEypj9ltYXKrmgpKWmXvc8m7KBQO73RYx+MfB/zXYLkQ4mN3G3B
Ji6Dj2QXlTib9ZoftLZEg9hPLAro6J9SpJ7no4nqxOvfe+2je+0c4dAh3pqY5c1YvRU81W9ZQxZ7
0YXGo02bikzS8Hbpws1uZDS5jTh1UZcENJ8MKBW5VuyYQCkmkhkPphY2uSgKfHb0Hm9rnHKsPp0G
i03WvLCbccBfVoh1+O2JAonkNdAe40628blyk+TECkhmmfaaoSTj+SakcyKxRkihQHCj+ctrkqBf
eRYIOPU5O2cQNJ2kbI3u9Ug7ITekRrx2j67FMAupBONZ0qERva96sJHPZ/br6p7U+1L3YfCF7QZO
rQWhHh7K6AWhfJl5oYIGUVqGKYQhasGdXTkVdfkOixyH53zdEJYTFAy2WG2d+l0qR69SmJLuIIU6
yuPQSbiLd5fa+N2CSnDW4C4sHipgyYJTWf3EdmUvQ6ioO3HgNdpG15MuY0i+T21EWUqjjjzA0px3
06w/xys4gNUNwz43RMQhOuGFRuXqiPt9VvOH9hxdr3x1GcjL0kmuuFkT3Qp8cg9NcwmNbndd1MlM
r6iTsHpMVHceGvGJl9VdYvcCYei48r9SSd9Dge9kHusbkVo4fIJXQz8jcaRP0DUMerIIk6CCa8Hh
OH0jlTGRQAFO5wXckX4fzN7m0ahP+w9gfKJ6PgCgaYTK4Lbzzlf8MxAPSGxf3sgMXbu4ZcU2/MGH
iFYFTWP1u1Z5EYdflsdyhD03xPLZwOnk0hFXwfifTDftEZO0HSAKzrC6PvfSG44mqkXpmGtXpfY+
zaPYhIP03QNqKtJHXld4LA9NSyEGnWr5jjkq6J/WaHcf5Dxid9HR0Gne86do1zd5hpveFqqIxWQY
0y35ad+vKWFdoAd8Jo2Dij6ac3Em16d/SrXWwaV7+9TEZE4fucqI0GPg4iulDad/1vthfRF341Dp
LAjlcBYLmtb8EBUBuJY6nvHH9/tuPshn0HvYJBLByWwqvnuJhhLNtoJoMlMFAL8nmvsdIg8/UFv5
agy2Ml/ARvTCD8Jeo1tkv4PdCvHSFUfuxCBQPhm5e4QoJusDECmKkLt5mw95BHhgZDf0xCNFpZqp
HfC+RVs5vbSuEztMJSe9gFtWg8X/phgOrdRXTbu0ZpuxaqxXH/EjQsC7jm6ODc7O7QRkO4OGo10r
1jK65RQu1SipBVP7MRXpL/10RBcjUskNyM2nXTb/hbi8gM6g9+a4D54tYii+AKuLV+miuqvC4EmU
TWQRguB28iZvZxYYMNdL2xXrB2/1pc7PxdUuYyIHg99vs8yQeKESuwjnUEPrmCdRXhkhB6seUsGL
YYFs9u7UxQ9ZDyaOLGBjH2gsNZeoep/UUumbheMc99fqaqYIbo2Bov4XZWMxDHYByQvc9laCjZqp
5CvzSnhrkggOUlQPe7FCEviEDoRgdxFbSqidhwhQwjhc8EvamGKLgqA/SopjEtJVRvwZoUtt41If
BaWjPK8t6pNB1btOfN2+eOWLJyhHQFNwJEkDiIgkBk4Cj+veY5JCT1pMtXUNLNcpMugM/2+fvjAt
Wf9JOjADmF6d9sNH74FjtarZhWUYkd+/WO5eF0jkohNlkOYu2lQJ2V5MzRSAZpZVhaKbds8UaaMs
/AGiRUXw2XG1R8Np6GrcmL0bqyYKEY30cR5AjFotogxqijy1cEQSzoAXSAqAIodO3M2bivLRgMmd
VZu5FLAFv9Bxu8JrAy7/vtvL6Qram6FZs8agyB8x+egkXY+cN8O4kXmLLkGpIeY4CcmkHeJm4dOs
1PRuIkgNsvpAjPF9nZXzYgJK1aOV2ZwtcH+7n+9q/utWkU4IBZ3cANubicFMZzwfNOT/LBqXdcQz
7uh1ch80aiyc5P40a/GwZKpPg53jRwpKJnxAn6EZ2tXgeiADrMAXN2KnVYT7+35GxOdH/YzhESdp
umL129G8hJMG2E+9xg3GYFan6K3nbhbkBREtqGzj98EPaFjFfESbJOcU0cnRDzbQ2ia0hxC/OzyO
z4IrpqPzeDT4P023ETb3zyv/qfrzeJG6XTsS48C3//GImn3OSbYoJykSSiKkKMhYMfbvKXfhUvXW
+3kXSjIGNefeKxjgEbn3oeALznSIl5Ob3jV6cV+s3C5ZYZvIBpFth4gBi5vdZb9pp12eN4N0iN/k
toM1iKVRNAQJeTTwKXO0cgT4zrD0gnl2gITyqcWrury0UOviJsmen8m2vLbqtRpyI0otAQ097qqP
t5u9r5+iyEuicnetITrRyTiOzzDpr2tba/kB0FMZMXj4TzUHR5+8I9/eAK0+quSisx4Rb/7wZtB0
FuaZpDO5rjarOw/NUtZROyRGXB430wSzudOaJ5kItHlIjzJ2Wfjm4XsNC+duyBf0THLtzZ8Oj1nG
y/bHC5Zt9AhaoocCAdaIugxB4FVXZ/3f94xZV5sxbkqtAfpH9RcUx5osk/vmb7jl80cZrmdJ01YD
hIMu0t9hVCKz69crD3RtWeUDo0b2vBzJNvcV/pBD2Mk5mVk5UPrSpG6buRfAzYppSRgEPxDVVSGv
m0Y4A9pM6TEvHmvzWAW8XTttRiB+zuW/XLCza8NAuTjqxTTd2403WYXSqfsFxhdtUd92S7z3BndW
un9M6hLNUuG/Tdvx93IWVrqOMd6x7fxi/Zq6KF5qNKUZ02FFRKBSliE2YWNprrG7kOt1zewcZnwL
Kt8zH27V2LJV+Kka6meDLFQFV2NKObdkaQxCNiy5dXVMFuJt06GebUNDlZRXC7oOIJ/W2jgF1ai8
zpfU+imGL7/hKZe8bUW1LIj8gS51y4tfatY7/T/J/gTywGFSMcfTJSVN0aNQ9AIgH4Hru/8zRCC5
DRk2k/8+m+cdLuRqgrEJgeeNeneuL4xVlbY7SoWhFSCwv9x1X9tQ0djXg2zkytt+zztmE30iC1+5
mUIa9WOYGdlSg7uFmQCCdkPvglHlroHH5WNqh2ISiQptwVgEK6n1BR2rH9I7bp0EZ0q2EbeHDsOS
BEBRoIz3/5MCHJFDCMcki1oKnPv1HXDYR5XmFC6h1eN6v1dKid8CfsqMwfHdasNVYdQn5zo7YxJU
6a2Q2TS9bM/QPTAsKuzVbkto3YiDRwymE3VXyu5vjzIQmzdgvRCeJ4qWhgsE4du7zYX14qTsTdC2
WNZOMIHCCWhDK2JScj2ZV8EeNGwzd+21kUiwa2DtF11o55QI1yQ/ldwOE849C1vByUglZjYGKcHj
iRqnnh3vLRT7D6BoQYq88fuI86aaGVoEG67WQ0ewVm5HV9BnnC/QxMV8DA4qWWfdkoE7/XDNv25W
22OVUloyYRdMf9mQTeFq/2HJFVaUuHs3L7txYJkj6KjIWrAtifjhBKNkPi88N0vJOb+6T2HOQUxE
04RicPNzTg+phC/KMh3QsGdUCCsKACuFynvuvwaua6ll1CLp0G/Bul6y97AkmvgFF0I+Folgtkcl
kYVi4Gotwsqm8k0esITZKUFSAHEe+IEeC9w+iK3f344ev5V+XcXH3Oesy3bzoY72FrOM7eN1NttY
HC+C0Bbbi2NUydI2SPHPFmBlfb6jFq6ckENDKA8aab0dp+SdD9orck9pgo3WCNyOLGfSC9RnNsuF
rNou4IZQsurPDnhucWUuak6a/FzKBEdPkyDndebTVu0ohUS4Wo8A8odntBg8a0kRXlsoiFP3eLIr
tYqghSWy0T4UejQslyaCyEIZw9Gpaq8dyM2LK8ckbnJZqQDC6G0dY1LBUGmhtVFvIG3WUfiK2Ena
kKnnDP4Lnh7NEJ5myZLS6PiBOlNZuAcyYdlZsW6qUqzPTf4QVnnsCBWVE2MKSM/VpzFGUSQREgq5
RNUEDEaXghTDXk7uYNKsCYg9XGvySCp4+D5PvpMxxnX7SOP6JfgF/vf5zk71WhOlaH0fnN/DaQ1U
4tw2e3RUesHjkKeuXD9wydK1aKej7CeMfhl1Dk+bkhXXOuvmBIVKfTqxblimvcPTAEYtbfduZiwp
EYLLoNmbaIXqgBm8QldBtAiDNLCrlm92DxM5KiQPnoh5su3GRAH+/evk3rxy8UQFDRpLJC5N2GXl
ucpqKT/JJ1rhmvwm/uoj1yGW57QXNVRnYIy0cL1f4xC/adnkWh7WDt+d/BOuUf5R31fqiHCZD0J6
p6bdhgy/uGqBsz1MhAHHxGBgHjR7DmxUS+iTcvndQ0AHg4RwXOF0wjnCOo/ziCVeaKUkRg/7MBjp
6KxhkVG/ppGAhF04WAB5anlvpW3rFrWV2XYO3nZpGA1CfYLmSCDjmELhnBsJEVEW9IGLS6WdyWR3
SN9tdEM3ZDCyQugPoyjYID0yqjnxNUaXrG76Wfk8a7sAKbxYX4HQTyd7Rda5nKDgDgZdPm21eIvx
dSBow+b6hRHQ4WRmz5+L/h9T9UJ5g1I/on10AU2hDmddA6Kq3izQxQzAP5wUzmKbGwZVOOfPW2Xm
lvDiH4HbgRLUC0yZmot22HuH02p7YUObLSUSqSUMp69dH78NR3y/sS2RRlTWWmUHo/jNvlUTn/SW
YYA0og11QwVPCfHRllwtkUMXGD09vYhJwjGe0tKoGoqOmokPg5nJ5tJraGukVvp0O9ZvF/Rghrxl
Nt6dughK5KjtavYmEFBGpbn2wuGg7nek8ezBiRSVbomTYm6ObFgKtFJSpAv07oBhMhQyL6ozlnFI
nHcCzsXNV9cTLGT7D3xU99yBsX/4n0Iphti96EFp34G/TcVSGbRMXk+esDxgLzu9S143zS+s5vxS
eTh1NtUBGwXSOUt+Yb35k9OckvSo8g3LAlvCIUUPu04m3e8NupB2IqhcFpBsRJq69JVZb+Is+/Dk
8MoN4pL6qdA1BfDyyQF3JrTiaN/cm+bka3WVj9HCR5pHJNB1OawMYeZOBW6UAsCSqMV/kKJ3slqx
Zht9UiE5e2tyqhktuAqE3fStKzhokc+StfM2Wq3YaGtPTV1EnUIPNRUCzXm81pLh53NFaD5HWqWS
CgCva6N1fFuIT5q279ULY8ZsV82+z6B0S+gejeGnJZDKN0Tx0ZRzh+jSkx8RWal2OYU+pkRdJDYw
HeBX+DjpD9NRtiYrxcFFE0w1Tt8qmLBrlpSOX/gvVtigIg25Ym/rxZ7wHmjdlbu+x3/I66lE87Hj
DNlTHEpV+0l2dFrW78aRh02Oe1FlCAid4jCyKXgSioKbiwAoS0deoBBG3dhIgIeYLCIfGddXdVLK
iFWHl/Y1dpoABj2ny4LcoBnQNi5p/kw/up3E0+LYEaCI4MnMBDCASd2q9YsMnwnp7QWTyq56vYT+
3+xoaRL/bNHM3q4mtnqXlATfeKFKXNit1Nxd22tX2rHPC9Y0XOGgyXjcHb8Uowiu3fvApnGz6FaO
lLC51ZJomfPzqKGnjaHurNYw1o2wwdJpD8I7IuXGmEC5kjRr/fy2JG2SA2N8F8i4kXBOIrkyv8JM
WY38U4imWBWVLfS+kxZPzsPddquthSwzpkAkDzMoICvb9ZuYpqF61Jr7ydA/fSuUTRBIJ7UteaLQ
bvCOlWDueU7xH+Ih2sgOV52zF5+hk0BFr06XpK4E3xcni+hEvrEpE9KzYa8dnyzjR5Ca5hzZg5e2
Bf4i3DKv7Ex4eaFaNvQr7qZnyZgDwmsjs464to2z2aJQozvTWPBbqO4/b0FBck028u7XFjC50Og3
M7g81UMLL7JrwNWyPZ/smt/2KvuNLJ+rqIzeEXrlOSRdAUCZX4kBTGykuzXnpJ3DwJ2aeKrjS2ss
Ojd5cip1rdD4d9TNix4pLXcErO3mhK4lA9bPEITWhP2OracpKN6BzLZAahL7sJX+/f5Mn8rjjphB
qNumTQL8G2DLe5pKVGndzu1Cnoih0UMZ6zAxYLskZnAQgIE7bxfE6Zx4aoairJ6hsVL/R0hSrwuH
AdKB/CmsVoHx4+NUiYpJcB+3uB2zipEmaiG8sKKOtpydeoiTlflfhjWj6Mu81DjCaxFoZPqtsEEg
2EcfSiZpgO3ZHeFQL7YRBXcAWgm6xzO7md5QId8ybkO+8Bf46IZimmw7Hb2RQPQWYOcAQD4cMcbh
EOH9f9OWVI9yTUcwSOnCyu2S8/0gRMUUbsy0TecxnptuDExr+6RIIwKf+JsBw+9pgoRxvB86GUMh
K8hrIvcvLxaBDelDyJMf2TSCDXoHPojwcdTYO1VImeNUFi/7KSG720dHEjlbSlBo8Ya/5v6k8kx1
wkrAFJF0AAasv9HkplGitp5GXQK8EGPTkBp1maKB+oCzPKEphuGjm6o0s/lOz6rcwMM0nS3iTcD8
c4PvqLWrkBPC/Nhp7/7ZAva9ifS+ir2jiqzrg36YDJfPDt3U2b19f8DufKLOXP4Bm+FQ1oziGSAd
mnO9CUw3j/oTUkBgLOJIe+DKwVGUA2/r7b3FaZ422zTHzsk8mrFPvrF2Q8ydJmdk6zwln8pdLya8
oF4jXOM8D7OhXnrHNdGMyVHvyzziED7sNKhpbY/Vd25tWAsdNJ+ZZte8iRp46pcRPuFo2RYcX+Mi
OaafGoGSMSgNTH9dpLMIJ5aNyi3Nh8W0XKOHlK8U7nj5vn6iACUzVQ+C29HLSXd/MSmoxyXzuora
TxxtkBZaZhTn6no3PvvC5W9yw6i2Q/wAAVUQWiev4GcfkJRfWAPY8AjMLYs2nJ9XjVy52SFvXpxT
NyfGoz2PXjtu0y/FEMakqh5JFLVWHiA1EDUm9zp+DEp+l4vMoulPvXIss8rLDERJI9GoXVFvccdw
QicKFHZSRGGFbbP8TUBHZHcVtTTdCs4olmQfLNYfdPOk2dNlozOzMZYa2TGCq04u9OVgmk27658Q
Wo+tZYAJ3HzcoOjfPogZiQ1Rfs02T5zr9g86rMkVXjivIeYA4l5MB0DY485cE6qrK8jiWQEPaazp
mMm8YT5o5d6bp/KAbNX/8WaYqlrUn8LDQbZsrU0mB+mTGcf7Saxjd5oipqyHe3Asa4DabdUKrXAK
02I6Mz/4bXUA2Rl9SRVpAC3jQt/jne/2a5BgpUxfHQVKDsRBPWcQ0sQeLmPNQDz5TpCYfGiZryNQ
Td7n5wfGor+gQhUTJJad6oPqlrEShNxk24qvb9T/eoofEZ0IwyIsxxefxJhs+Xpfu7Ru4x05wA7N
iRjzSNmQ5htZYvuv6uJI2cILWAFs7xzB109NTbHigJzCA1IffPzCUKlyo5++kZ+MnghKy8SnddCi
YtWJFoQm0nsQkt3CDzvq8FrARBC2LlbpAIcDS+s+SZpXiILaZfxnUYwXn+tMVIyeAhOA2RavHUte
Og0/+lHqXq4JMrZJ8huYwxthfXHZuqKnZRV1BRQj7e83uRnELP711UtFaMIxJe1GG56rNGi8ESRR
5EpkgFxft6jCwtFBvScKKIRAqohumQiFsbBHhUPchnZ1m5du0rEkUVRvMPiNTrQ3cptYPA7m8pmx
wns32yv69nFmSn/q9X5NR6U5clVGk5mGQzE5iGBRLw6Qe5IljnSqeGe3xFap64zpGEwYasIbjfkt
qpoRpRT+NqsShVJbX+HTwHv14PqlJGLbhUW3LXpYQhgsi0QIZOyIgthXEDblU1Q4ztyjiwpih1Xz
AIkfWi+mEHtgFapqzxVUL6Dk7ZuXb32QaG/RGeutXhwSiV9idSJThJm+2YihqDB7lOmClAM5+OVl
PGiGYklugxA91JJaXT5lzlvxgxfArlkK3zMATrCxV9zsRLefY2/33SCih+3rVo0UmU+ppFM87VmD
5eXyTS9YZra3FW2IpZZgtql6CprQZBG9x6ZiiU5Semk5dBMOF6em1si53eTSffsE5L96ispLPJGx
zCnOy7K3am14ks4hADFglvJr5eu693+VTvFFIuU3RWlvVEDiB0z0xLrLL3TM7a8QYbqLHy8tiizV
dRlKbQTBsYE4FZjjzi+pDZ1lNe2TWp/s+E7dgH/YjOSq3HbAF0MZC1FwHk0ratsQ/AccktwUd3Vs
5OTsn1JtTNydquyw7l9r2GEiEZPwnUFI+I13A949Um0Q7kVsLRaLJ3ZSnCdTg15HP0TeK9TAcwT6
v1hYkTKf0VSndZ3MjjhrMYBKCWPNrSCs1RIDrviktiwUDLp8iOVsRAmRw42rdpBREEPICDmZXhJw
ZY6ePz/B6HoctgkbrB/RjyIwbRi2XdPFW6td+HIVaXf+ydYh4FmqZDJnMIGgyHxvU8vI2Yt8uqk1
XRp+IaONNSHz1ZbMeatt6uwKG7wI7qL9IpTrE6w+qE9GhGVRWf0olFmnNP9fRPbeeAbU5PgF3EF8
yiEyxlruQMujtArN/YuK9P9D8trvz9Q3Z5S6dv4U9FtoKX3BCEeBQnsKEBA5NpDHOZnZL/8aYxaR
XCc1D9QUnTLHAHjg8mU5EmWbYtjAiADcll8kHwWzk1IQRX4n5aPgrGqRrfrAgZ5bYA7/x7e7Pk84
Gmulf5QVWonDFB5PbwkyEWWekuHij6CDzTufz6DOTftAUyVvIGbRwgsFICi6zch8oTlP7+ycz8t0
`protect end_protected
