`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ikj93e9A4VLdlzvIk0rVX/rEjKPQTa3gVlC0+sZtXPKSZcMmqk7Di5XEs4hnsMV0h2+euwi9TV8d
qv5g/jV/1Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ULBoQZamxgCvSlaaHpFPnePWCi0tAWiHDHgXkcKTObIDQGYVuKt9uloLAo9889JZcYlic2hmqFWP
awZXXoC54Z2wvZL9Q8e6aKrcEOQQ2Famv4Mj0iJE1pyxVjvwbQuHM94bvltE6SumK90zeL5gvPpx
UokcFz4XxSJpYKi5gGY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZLjtAn1Hez2iZHvCg4LqFhmlYj4Pp/ljZZ5odgumpUDxQkNDff0WWcB2NNVXZMORoMaw9VOBGYBA
WRvYEFRZ4uNSN7SC3HOnEHo8Totlf7BdgccVKH4q1NL10E7jS/M3JYBHtL2vK2124JbR8ROQ2U2Y
ySuAc5ik9yuLCXGihkzBqpJiWwgiiA9t9xW+0aw98h9hjuaw4ydli/Z1eiYN6Ec0/kFEkRvUAXre
8ByPErsFGq8LonI6ogo9J2jrwai/J71tIDaulVWavidy+ojyxXh+jvS6ABPlwh2dUcJOMkXCfyda
+VXn/hkZs7q9cQxAzHJWUiIaGY7V1+V10W1Q9w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tNvmI93w3vSlIcuPIsU4KadFeYlXFwIsGx9WIbhGOa6ttVl20oG9SxSu+rhXXqAIO29/QHrb6lBn
8IQ6dXSa73vuOImlBhoswOesIfm+YqZ/YuCR+leqphdPn06OW6xPgj0x3krWp+OWSF/qUspCpiHS
dx1WYyVUFt57wce4nKw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hjnbO+hchdNL/mLdninO/RoKMyD8zMlmtwFSSN+OXunyBXDW0SDttglWh70c+77QsOty+qGYAj+1
40wtW9PVxIpu2XR24Fto772krn7gYBmb28SjNGnUMNpDHutw76ZuXd1RiA0JJrz83oCvmBFs8OjP
qS7BHBNnPkdG38Smbz52pHNcJ+i5Wu0IvT89DRbNQ8A1WjDaX6dDj9X7ZubLb0rOEvA8EFMKrIib
2+n/Paw5/ff57Ipi0x654n8ywQ+QDLn57YtA5E9lYRtn76mvEoEogjeUB8fipCjyGRKTcojtiAp9
mTa/LLWL9+m10t5LPlhgsesTZtYGOAcnFGRstA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11968)
`protect data_block
7T59uFdk9Da52VY2RqMBAHrQLJpLzK0AoifehJybaRoFxGXAi/Xfb+/V/qyUuGAmzOpX8uKiSofn
3Ly6GC5nSHhLxYvDSB1pLE3AUyl1QjhP7tRPalIQfmvmTNeZiP1zn4hfunobzjeXWLml3VxzuqMt
/4TeJgaQPZzlsDTt82NhMHbFxV8Q0Is/5NQVGqEexTLM4WWjfyULXOqDyu9dzIVJ7BnXXQOgyIU/
ClIij9OSnpi/bD69uoACgnKUGb3n0YLp31ez7M92ysyVk6P/N5/zPetJrv6UT3RlXbV03HKVuolt
ev/TQ2NCrzygBTV38bIO5Yahd4T88F8wrgbpKW/3vFRd1OnL8sJO4Duyg8nywluXjOn8ewZ8Cyn9
3E7zw7cuIdo8mhDITGvO5gJGSRAJdnhSSArv7G41hNPt76651ig5r/NjjIMvly3itXdXXMD4tTMw
2aZJe1DZL7uj0WZ5wNSmMyvc21wvPr+q2v4kE7a9qtvxXVT7EgOLgU+6e0lsXf0gGbSiDTXV4rFa
1GdRKhCaSdOdcxgdSBtmBSGA3nq1aJOqBXQRRfFXJCMg2r4t3Pxsjz3Lk+OjuXH2aUCDMW7ZTZBl
4dou+fneAStlX096gyMDZO6PIn9VyO+F39lT0apmZhC3EaIIn09ymjZJ1vMBf7ci+aav84DbiquW
5z2MMfw3ofyV9I7hUrdqu/ia6XOmqxnfZzlGtNDhTI5BN5PFsa2Cfk+i3P+78Tg1TGvmUimkLcHP
/C4UWJlGd/tMmDmPbqp7oAfhPpSulnaUfuWCpfHBrhkkAjzoxQuZuu0sKS8qtbYkRq4mnztF+Xz+
C+ShZ7o1k1ORgC+szwe8pi/T3mjzerCqBdNbzQj9QZ2FThud6D7Mnrox9YIZUe3/wlBQ+v8SUou2
PIZSX3n9jiaVqrgwZje+iuRtzz1bbLstaMOHMBDGLUIXzmu9XCmQ0Yi1aXxId3RE2Rl/xVK70SQ7
OVHPKJNUh8cGDzaZN62+iJqkzseH0lfxDYY0DdJzgMhrXMZOF4hfN0aFrxcV2nmtB1WkmSJOzTW2
0LNYoQ0M7w40RwOYSc/+abPhCnZrdpCy3VYf4iHQkXLJ2LirTGnMjIoGdDMwgtMLWpp/VZMkwn0n
THV2d96Kcy2BGR004YxZ/jo8B7398B37KNsLPhIa3LLi7406FyAgOe2yVcMvhMSdlca4BSKQIiiF
FGo+IUZnN0SVVh7Am/Vui5l/wXFGHQZ5jRFSxUh1+PdbeFa38M9BGsHphNvAa51J7QnmQlcYfoYd
TShCPnLYkm8Ma74emFola9PLVPdjhW/E3S7oxc1pDX3/nC/i3IJ7D0NYheXktWCQThSa3sgIhi4U
QGbRAmWp4C5rFHa5D4AvMwnuGc0Fn5hwRD+vG3fRzPVGEXHNvMZf+i6bptcYgpRaDjGlvCVMNr1O
gTux8HRojQ+1k/C3IVStLkgykZ3EG4B6VArcNz4tEikK5ANFvkqa9UVILyJh22vS3AbmvcQbJYby
Rtf5EH+t5jro7UzRT+feql1DPT6PukCZJMWjdRWG0BV6eMPQRk8bDM1jQ8shxlaoQCpPmy9CN7RZ
AkdTUtaYOn5kzDyjnKJS98l85/oRnRTzKVAln49tH8JCI+o1Hw1aCHy9wgu1lGqEl1lZQzlEDRPg
msZfLgD0++Dq1EEqovCDLOwEg4vYd5WMo59fYe9WknA/ifP2eLewkhLtri8Cgk3J2BKhBmtgcZsY
PBYQ7G9mTLcgaRjtJm9lnonXHjjEuD3Xf1RN5+e7FdBgv86TguTt6RUsqAoWEvhZec0qPYa1GZIa
TUQuHs9AX88ajVx+/08mLJjUofSo7pjbl/QhjwOwM/n6LoyrJ6cDTLHXU06MIBNDNuBfWBDUpChn
0VH7aWRalGDlFmGWl3SaIdT6APHBHBap9WRDWs4zpAwi0XFgLiqQtkU578mQnnG6HepanuUso4bG
geyaQec5OUQ2v5z0z+IK5B4KiZXjdvKtHJmSUfbdI+cHgbxvMCzW6zqMNbMlMO2sCYw5rTDD7cb8
yOCBgPKDfH2AUoQ27wMW1rv/LohkJwgQVYeMHMGuJC3BOBQ3CFONMRm2g35opbNp4N8zERTnPXCG
nqmJRvQeg7hYlNQdH8l7yFFhSDbpONDmaycQ+4vstmRZgjG6f9UWzyh3wLpt1qWd3EA56xtWT0QI
veYW/qxZ/njk/1ILul3wWKD9YDiF7iU+dCIs4t6a5A2bZ14qTQVGlna0VnFNqylRrvUrqwn7Glyb
k38dUbnJ9YJ2OU7ujU2MTsnMviam6uqbjHxvYC8j3TCL6HzQaNCRZ3stVNSXlaNJuhontXP8PG79
89LOTdKSScjfYMdR3DbumyDr/9ZH9vCAHkCXdBhnlquiuYB+4EarE3oGV/lxC2unmnf00uquF1Xq
g6C5YVM68yV2jeDxZYekuDqvd3/aHR75WZFGJcacBLVBwqRHBqS2ubis9U65El5N4NcNRsELTUSZ
GqJDxOdAFeIlb6DLMh2PgdMo3vUNZFEf0G6zM/N/J5+vhQTK4quE7tgTpwTOVzk1JNGcW1vPcudN
8JElMChpWs81RX+5x9V6SRoVatyp87lnGOFH6vSC1wqb4s4bPKQwmFPvQS7SOBR7Boj+iIJ4vjPB
Jf6c0fusa/IoYORKXVLjxYSO/ZlozapSxOkvmW22xGG0Rj/SyK2Mv6DFg4WoEV/G1nXR3LTyizbj
QL+uc3uTSEGfdTuxT6i+skqh5W5bWYWaLHE0Lf5vccs62JG/V/T5SY9Yai95eMJ4SSP1pdBoFXes
7CtacNYNHgQtrefMBFc/Z47C5iIgVPiaIPqH2o15vRvqDcgp0o9BMUIrbF3sXj/PKMLUMgVp6t+v
wKgY59PXRBw84iTxG/6X0Xtdjlmk4K6f7zgkRs/aUDaV0IkqIfOVIATBbzkR5sN+JYCN/b7VFeJc
01Hz1X871B9dYGy1cyS03tpDv8klneokReUF1QTKuByLEcXR1LYyYbHfSGExlQtas7N5qtTuqsP+
yYaZP3emIVcQDfIt/r9irnheH1fauqCIgI+vXg9hg3ZKUizdVyAeLJoWm9w0YuKRxeUWZ6pNpG+2
7eId6bq6HEs+mr0vazfkLpQlIVPwcIlQhtJ4PTmX8a42vvUugTcBDrqU6RoocVRGOTyZ1aAay53x
mi0bnklfjYfLSGiKrFSFfwQ+HvSf2r4YIlnwsnOrb1SIwoYSG9sNQRoikJ+39mT8gyAcbhFX7/6A
3wHJCb24tmb1x7GlgbCAkptMlRN88dsKzTL7e+R6jycEiY7puVKYXqLTpTvJoDIr63a45ljE+9I5
beNAyhlAIQNGsZp/JyGF3bgwSjMJeAUVkE17QsVXwPz5ShyohGA0a/GXtKQ15VqCDBed4qR2vm1G
Cp3B/KbEa2sZ/41bxFKJ+9pMXVIPORbpskedA3MEak6W88xFZBVtRaQAqFAYOPuco0Zk9mnnAFp4
vXaopBw8idQ9eGkcMXFGrr5Y9u3al51/NUc9sVOCOA985eLh9kEQSdnavm3F09grqx7EvLU2NR4L
dx3wa0Y/raalRkCZnV5OHdGDo0pL5S6mJuI0H6Z4NzQcSmUYIYDBVtB6TxINwt8lv6Klf04Aqyzm
yUQFluiO+PE22d4olEpYnwk7b0GSm9FsIs+W+FatnczHaKoM8aCJn9XJ+xM8aVn4T8dv15SMGTSV
caTKRaCNbK4IXqX/URO2TQqM+Yg4PmFw/v5zZQIC4dKZGxVaZNyJs7ntRF2sWfzI+nulGG/Qksvq
kQOEwbRdKjUox2joqM5v9HCaUjLSd5vsSfp3eL9YrFFejqlDWqkWOEGSnSvQseQje0ZtVKUaxM0U
EVp4PDV5bdRIxiJsPBeWTdvPQhQ7ldQ4F7teYqlY5bG3tHxm0gu4GgAW4vT+CXHhZPt1Zd4JbQVQ
u6nOIOHGZ4wH3UYQzNL0choREXI6cmUaE09yE1V5lSjCu0YO0laPjfWwpaVPzB9HUy67Eq0LN2zB
3xAazlW8tbD99OMyJOeBCrfC+vdo/m2WjpmZ7Keq8kJYljpYhXo9VYvb5CJLdG0tTQqBSsKDOZfj
MYTeK6kJvYgHBU3f7d3cWuINzXePBYRUMvtFXSwgxTFzD06uae3toknT9ci5QUdVNd20IZDxME9G
f432H+HZVmrR1gcG0m0X8ylTkvHHH8TADl42wLGeT/P9xoFFg7jyPodHtNHboZapc3c45sTnhmPW
BXAI/TCh2y19uHRBpF9aZrAK+KLNdJ7VMApq9wb2p7TPxwKcF94m2Njh3duKL4QMFG2htXnGHcl2
gkuuR1tABrEkWWic18HU0aJ/geXzm/LmOTOZ+clq9Q1vfiT+u2EhRVv5ThuCjL1CmO23kpc1xBSc
lPppW3+AW2D7DY8GrhE1A609C3rUMq1RFLZvWY8N0afvtFHhAaTA5t+6WKFLGcgwoc95hgpGdBvM
aKwUrBkLtthvczyYMWg8LuIK2q4nUL9xaGIQCiPQfsn+wW33RcUx+01Ixz8AQWdqwJ8Mhxo2BJxh
tj6mCE4ELNaUntuQn5BXz6gupDAWLn3L3sRP/ZZBF5uewYqhj8qmYpwr+KeComTxwuANbqM2458n
IEUALZr0OMxs1EjbzoMXI6PkO2aJi3Gaa3qTCZCNzc146vQK92n/JURWgytmulBY6lDSOzbcxG1b
iH2txLQmgQfCAeHqpD+dX3gS+44psfNO20KVIv52MYyQaTC3tqnG5oNow+MxIYSHS+I5JSMKpEte
V5boTfg9S0nBZVBseQSr7RJ+0cPQUNg+61iJ0segnLDlD/R/xKFLKIlQSTNOJNokmdLKl/dV0Aut
rOPREJoYemwILJLoUPHFrMmRrSp87uTPHVGIFPvWoNCQoOkr9G49/iaWxqdBk/Lr8sxKr5cQUDXA
eQ9h2EWe7rQP3u58IQim0Y2CLxdCr8m5lhCKCxXcOuHKQukBsBJKYvQtEVf/+sZwT9D7W/loUjDk
DuOqttFBBJqd+8zV/fQO7lVKHdJhXrG8+Jbm0TbYALkRQnkwxxWbjsoSvsUJhZzLh2aFHVBrIvXg
Ryw56HMGZN+o6VsS2iNInsykyemw6bm4hkgKUiIdffE6J4kNCcYhij4NSXPq174zhUsQp/hmr+Ye
D+VXso9Hv5e5SkDKrY1wj4mQV2xDx2RFuDuv3kueMpKJL123cmgqp4pOSguurrxq3u5BJJNNWwHW
6QQ68VOmMZ568gRPcVV2AZWQo64fia22ZRyMjvytc+S5uID0p2s7VKx80LSD6wV0LO524BLdClUT
3rVoZwT2Yhf5QtqA15aTLj3vIvLLsqo+DaxpYe75SjLzv2DbI42KY2CQ7K5AawMHFTUMYVSp5PbB
vr0aRKkupWLHZPcRCXGnxyBKTOmdPD6DmHOyha/RB+hgqpUxghLbifioeAxPnWtUrxxsAAMaIdX5
I2WMeRpZzjqyounmxOfI2S/9/6bcUdClWdM/vW6v1mPrc5LPQw1zgKanu56Yv9Wl7YtaeZkT64eq
2E1my1NJEOYUp+wWzyk+kwp/adElX99teTf6RDs+zyWDZakXpsOdxaxh4P0dJ5ngvfcIl4EoHtB3
ObEv5Eg7Vc/sSif/vlrdUTeJ02/t+SuphHkDZHzXYE9UMzfbk/7ISKDExeVmDTpG9C2AoMv83FkH
eXPH2hkrz4Xo0z/rFT0R4Dffx4TUvnSsTDblVgePtbeE7yYLg8t2gKmezWzHo6nrZXZ+fFVG72Mc
JWVFfemP4+TKGo5dxaz0ABf6dZ3qEkSRPu7DTkN7te/2/Zh33CxfNIassoOwItvTxkz/p38CErJg
5xwozoCFgOupvFOeS0DVyCAR+H/PwkpbfPdZakBCKLfXr6h+j6bZAvXq3Q05Dzze6MKuKXmIc+lq
mV1xB7guvNqeN6n6CVq8IjhJoDxpITvf0pwgw6C8+fzvQQFkBN+RKbd1TBObo90AvqIGYZ/KyiXL
dPcWq5BUcIK/i5FBhIq9Dksmew/jeLdFJlpYEeIVs5HfioYbchwu4Nt+4wKJiBQZZ4vadDIXsAg3
kKz4oauRpdr/JzOlz0h4p67Xc4x2Ku949oNFbV3J70CVsGpIpRJ/rW32pHds9SwYhjNFt5dB0udV
8wfdXAvb3s8YeDcSKcRQxfVfSAyH01o1sj0AmXCVrZBYtWFPLqczmPMkgSbhgHLkT4pH4xT5plz7
Nz1eJzSEE1qOpCrrj3yMELC0Mr04R//SxiH5I5nkcaz73AB6Un9Ap/qKXU8GQiOl+bgzdP8/Thni
kYdBu97G+KZS2bxqEWfbL63eVDF2d38qmcXD1VRfehovKThRcndN/aKVBKtudgQ2cnp83Qz+KFI0
32B84XN40BO76LrsNJkezyXBgeqxu8WShYUH9pgDax4mqB7BRE+qex076nK8EC2uW/ENZxqpVFZV
A3/kMdVsNPh0cRGbLFScS1Cr5qIlK4Fz6hQT+/r2QMzSNL/KdpQjB+3Hzw/7iF5rDGEVoRn73Gm1
UxT7EQBR2rToRQogwhsdD+EFjaIeIvJtLXCym0Piigc3+HlO8Ate9gP5qiirk05eFiiu4hxG1hKW
P555c4fS5SPzdwB95pyyR/RvGgDgrRcR3tHumCbOkythDGx1vOl+JQB6POU0wyVgmJGZxAMpusDS
I0UgoM58649GTJCkJJkLTA6tdoXCslKZ+HFLYA0YySd1NgvJyPmXE+PB372bpurZkgB553hyHiYz
yj2gJGiVcXdu+xiP+aKp4qVt1slL0p8Wukl/wlJKwc/g+lfaGE/q/Sn6DINYZEryEZzbatq911kk
MLzUEX0S/PmEQaZV85pmmvSx/EDAEV2TIe0QEKjXb0CgT5BIctuytrU87spcMD6SxfVf5K1dPlFq
jUFVnIvElz0xeuUwMO++DIB/uO/AM2gbNzoNtlpXr2Grt1R2uyGbuBcz6QVKlN9tRokioYJRLWpv
OeDSt/GGI0NS7m162VoOLhvEdCyEwfyoiKHjh/3B1r9S9c/4op6Um6uMzDeJP/qnvT1Ae+AOaUlo
L2ZfLuIm15QY4y6bcnVkr/ZNYqL+gbPBbgKYILstLKIV31NKD79NV7PcQMK/IpMkpSYBF1LO/3cv
Psx1Y3+y7OWcpPDRbDeJpnwWe0Y/W4HKZejjsEMVGqRhR2qDtFslCIOLBZgUl70GAP82zg/s1vdq
P/l0Z3KviRvCN6w5scqW4aH5AFN+OXTRdjW4VKrcC0haypL6Tl+xfADEKnNgwWKUmW8VZkh0eg7D
KZJKp0eFYfTg5hsEe/w5Ku/ofLMbG7mD6L0nnIwHQpN+r3+843AK22tQcyXnxh8eW0OIs7lW3Css
tG6O6nlu/S0j6HTJSkWW0VBVVv59crFHJ4nKQX0o8mjlWMboNNyTfbefa/3i+ykDjfkY0sZ1vQj6
jyN8oOd8lXzMmiiLGYpxbiD/qHRb/2V59urqMW7l5bRflvqsZmngggma18uhWKZG3wdL2WicdK5P
9t//D5hI/gLFt0Fcmcrev5kzmJG1/wpUtiw8VOvMXkmLyTu5s29zr5aJvV8IYL+7kHkn7MCx66P2
959LJHDh3HDZma1vHuwQ7k0n+/iZsiPCFj6uAe/r7YZPkdi6k79KzgPzEgVlsJ77idM0HPZPY7L1
mfMD/7ru4ozzfGkvEgBjgmmRXIC2aFDQ3DX3wamovGz0GFuJNS+ZeQFMMqRlCtFI+l/B/aFJyc4S
AxhMkPV8u2JZ7hNcaBM+yeJi9898phukUwCyoa81CPgNFEuegha/01Z1+KamQUEUbhXXhTFphlII
Z+s1c28/TrgduVbGVleXAKlawQJELjKQbqOKK9Ds9AaD3sPbDn+hmkGG7Unp13D8ufeuiRpPW1CK
zmkixMM7CKevs3qV0c/wTvgJXVS/nUFvZoVpe93ZQZWl48vv14tvsxhWbqf4pl2QLzMQj6ktANUT
BXogWAVrh9q0tHtwYQfgzrt0YUilrWCcEKL3yvQua1JCYLKYPhEapIx9T6/0ahEmiTq/b9m8egD8
dvvSgVYAwOIMPcXwDUr4+BUzVIucECTwGosRD9XoGMgDfHlcJe9lgWqpZqd21Osl1V65XKUlF9tc
/nNAaCKfthPkS4Q01/SQitBOvV7afvG7c5CyGnTJEbBhKzIyIlwQ3RndrKwKAezYOn0UL4a42dfV
XYb7pBfEygbf46HV4M+dwijez3q43SslexyLqohY7l9KlOxmgldGEzAIaDBC6PHP4oipBng2HmyO
XcnTPzxC+LrToy/Sr9WIRj/9MCJuCGWu7MtTi0BKjXvdIxxoDldnhcxPJI39wLI8EFk+CHaPs1om
uuXwo0X2OIH8xWX2a3KMc9TD9ozhmRIK80GDK3RbWqczVVfQ7jp4dZnR3QPKUMvzefuO0n6ePa/8
LMmwNx1ihb2+CKJQ3+RsBv9UxsLgj2qByrVgAnShb41nKo4K2g0hpj8cy5hRUAY7cOdKO1SWhSgF
XRSO6wcz0hTc9UeEw/Q536JczuoDIp3NJBkVLUNa6vvClgo/SkZoJb5vh5d49poiPEjbU7U7rdXl
BgfiiV+SS47viHzOPNhWdC34R++bzq51ZSHIodgC4XWK6AXHIoiCPhOwI5fQPCZGr5R89ADyN5WL
zWW562G92Eb2hFbhwdwBUXeKlbpV6bK7QMwAZzX3Y/2vTbU6cYpeHz2ouU3i4Wikhghe/LMbE4BO
9DP1qxRy1zH76BU/XYLCzCOmBBa7lG07FvTXeb2p1viuCIrt3wmG0w8AmbyGbDUhjC+c4JJGa5Kp
nqxbEDgD3ESiHasmbg6G6PBABv6WSIOpdORGGooclKGQ2SuF04FCASIiNVuWuIQyPHU3Y9+3xzeN
r2ZBSLFT7aGO5TGjGC7zc3M8YfUEz6uega7aikTGzffvNKOHznXCyaIj4/ZAnrLpalgDyBd26uqF
SPCb990vfj54kTDZGI8iPlLEnUgYpZOSWMI3L33aFWG6lucsZyMoEvVNiLAqtht0f10Z6x/7bN8L
t348hGM1BhXR7ga3t4ZGbTFPBqd6wTU8ofBe4xThH0PDN31otH/KOjSmYZHKk3ydCoq+F6tpEARj
EgZkggHF6yS/fFrKA1dqMWu7sejVd5GE7mz496h9+R2Lu4Gbu984WZ+UszNDqBqOUjS+8Ls1ItTm
IzcPJZvk7lhjbF0SUj5yeJSyD34nT0ev+mBjd64J4D82Zwngl12PDAO9TGwgdBE3teWxtFNFc4AR
hGCwjOZ6LYZq7OoVy9ykrYsdLOch5dIBM5VItqO4/l6vHckJEpTRKHNswt7rKO5fhJ217EGflro8
XjcqQpX/YahnlW6+hdEBsL2sVhGWrtEPmJs1eyGiHB2DE0eKoHGxdVAkVYBSHKj1OqvVSVDfnZ94
lfM1DjvEzdrEpwvScP9DI/pwII6c8hPG3wVRcgctjQW8mKljPpxWC9Lckq8pDGpcp1u6x3UDHg+u
x0dRN6dZ5gBOnp+CBammD1+MEyfsQYyrmcaPQusXmeI54codlYNMH5tfE7WOfZ1HSbiSQ5IuRIiK
MMF/O7zFmygwG76Cf1pn1A3qGCZsGLYkhAizpLb5L2gEWxTYxClvWpCUAIr+QDWizM2j0R789PGs
a3Jm7kOqcmiFEbvEtqflWpk6cZNznDt9kgn6NpRiY2SR0oEO0pWWxhO2JxmLQRT0zQleSsct9Xr+
rp7LTuKRAPYUYmawBXZOtbgJHpJijzwdSF7BdqM3lpc4C4TpIUJB2chbATg8m7z1zjyiAMJ60FOb
4tV0MzsKQqLKj9EP5cpugbCK1tzVA0FQ+UzdIr+HPUkg1OqobrE4EBEXOj/c4JBsQe8h8A6c2W0K
XRa2bXOFJgPnh5mEKIB9ucWGZ4r12KFktVXLywU7F0DvHly+vysCVoy8F/1ietDzsQwAFbbUeqBz
r834FMR68+dmFatmJBKWxXFRcClY4P4l1lN0z2sf3KT5UmSgT8OxHWgcQL6D6aEBL2z4ZGWamizO
5WfMcB/9RzvQMn95tAzsHQ4QO+8UN05/jFKeu4EVzrLUKDUD1/7tOZtH+Ymk2KEA9rwdQCJyVnE4
ZAWCtLi1slnEqc+wAEi9ceNj+X0NRBzvqSbdX9WYXuMbW2Aq9MhL3RHiKGlirXZ1dPorlTzP8T4e
B+xKXYRy9M8HoP41hl9Sm4tci4ds69w2Xa71ZEejDcf2vtGGIe9629awxmPywn0Ipf7+qtvEf1hJ
UL6RVFHTxA4vU8QiMGAwYqa2CpGUox+dX4G/vHAeOX8MluVfWH+qUNSGf52ouK06hjbS+GBm23wo
/POngTGi3MxucupTQcxpnuEopBb96bfBJNqm1F48oHQg7f0XiJc85WbpIsukeTRFuBOzbKkpUGko
CEayJhzYLaZ4N8rw4C/pZWPa5+qxQl8bOzBIP1PN2wQYo8m9sJSVUbV3DNmMgiNnYuEkksqxMD/z
mI310qnEbVj9jjKic3HMK/0KgJL5siVhtYoZMno7NSDFaqepf84VqprwZvOINmUriFX5o1h3GxW9
SuO/IU7kMDSUOXJfdMrk+XiMUn9tDgrtAo4QsluOPyDNQhfjySbhEx11FcQ0dW39taZ6aieZso65
kooGfkCjg7EYzlbYEKD+4fuxP3vGOUUEg2/vJoDeIhU3jfB8EpAycEovLwRk3LuyI7r0646H+y82
Ch9fC+gYRkCCOfv/gXYuO5Cc8VM6RHEtemJOTwSLOsSqnwxO0DoKTxIauvFGlKvX2k4aUezO3x8P
WcmZDuRa01bcx79TNQdkF7iXY4YbeBEJbUzAAIVbotBnyJDHhlcf6rsdCOl3qqnnmLm2/dWMLHKT
Sg7hv+q81zzKhoV+TfvAYCqQBMxkiCXisVaJyRgbblqSued7Wb3aFcSizAP5lUjUnDBaagY20wB7
ioMe7FnzGD+tBe1dnYBiJ30xU8/1Ga3ZO+sXfwAlRUVK7S2LZt4I7cvLCDYk4agUbH+j7ryj0C+c
+UlDIzEgTGj5MCoAdGpQ4HALQpSHqpu9bE9KBWqdldKydL2PaK7jbNrRl7W/bkPSNcJtVYSSsMwX
tI1ILmuzPq15b7cFzE5X/zLSTkVt8NbKdmrD/tWYOLqQJSJ3N05xtsp3wUfHlne/aTID9cunjXMy
oyQWH/0BzLVdfTXmEhPkYcHKXWwxITrMLxmxRGpB70wXGTkMQhJuEiUEDMFJN1FPR17m8QxefqJm
ezoaO97RriGut6bJ7OxJzxAEGCI9qA3jHxljOsVUUkJCrptSKm5GjToOxUYalboWM2FAsIq+Pd7o
Ebxa5jOPdfgvEweTwS26lsG/7uYfTSuKA4jpofXBUa2cd74FgyjgNCI2ufpgWAWqmzQ16jhzCfqr
a3K5gZpfUXqVrpJPO17LV0AfYt5glGUaS71ymCg+639UgMDdYTvOGI9b43C4J1CazVVwR595kfPu
yZ5hzEOPwYQiaN/oaAbwbE4zHToq4w+fATzANQTNH8hl5avelmsQv4zxtqqx54uAK13bArapGY9j
yDoCs391sNKiXaLwzi7eqO1zAh9jOJt9DxCe/hnuXXgoY8K/xWkmsH7dzlMi5uwOzRaNx6HolDr/
60Ky+Sc9pY5pRnGBhaZChnSrkN/U9VDqlUvzKbby+rHo2FB+0H7svEH9vs4V2xe3A5935CktCeXa
oNrgWwUCq6F8fBC/OjyD+Rh7pHACXw4dsrWn6awxqLCHPX9eglK8vT8CBH0Uk/3n3YetClAJRL0s
qDSzoRAPYF/XzVFJOtwhnO9pGSSmIP5ogIbnPUZbumipl5EwUIztjuf8wZMrx0B0tjR4L4HMDm94
V2MwvzWKNgLKgsH0UT+bxsmiIeM6OoIdwFZBjkhCCijPS1a2sYbBBOdxmyqVd4Uvvo/d5phX8KbU
TA5S25+IHFHDH5PsFvPnDWIeEQPn/aEQpxbxSy+SMI4tdS0XiBWdWIt2LrS+WaM0rrBfYR91bSr+
AFCw+76aoq2r0JMqLVQXGGgYIx0H7Df4aRgZj+aImQJPiniRjNjufEHYO6Sw/ul+fM2Eo3tvqTK0
QDj4gdzAnGduD6SDadslVywJzsa0bRfBXKz2qQScacmfbUaFK3sX8hM4FLuRGmNPeBSaAavK+YKm
bDAsZWJ/OmsaMBtT7A2scXz57SE/6ss43bIT+rKxRpvzhcuoZqmUeLJ4X0YFahWwqSXIMlU1GwWU
r1+n4ZlRpOei7amZ0l5OVrDX6zPAnRn0C6x4Sl8zHbyLw1dMLTi0qJD228jKsiEpvhraQSwuihKt
tc4dY2cPGB5NyJ4xIHMKTcDWFi5Kg361c1gfHxy/UhoxW17FC+1f7yzotyDrPke5Fxq3l6toyxp/
pDbhY+RHzTnt1VSh+YRc1Q9m7eBqd3wvfxf1RfJOV1xP8th+trrk961WkPRrgo5RiHQvXSt3RS2+
ibVMD7W90LdAYlqEbGa2nGFQlDUgV4ZY19tfMdfw/rPvx9sbI4CsqPANPRSer3D/bh3PmtIdC7NZ
CdFmFvQS2z9qgvDLywDpAN4mIJEcVXDMF4SQ07dbc5rG53+/jdV4/SZ86Ji8Zn+BfeGgrsPH7Pp3
jS39YIaTzSeea0xddg9qTjaiepLbKsLTkzm4f+LCAcdWZMSRNMnC5ij02djbdWxpRs9IoofThqYG
ErA2Nwz1NkAyf6yO1LnUFg7LYuidPwUrrUnW2ddQbLemLDM5oAKOcfgDaD+SlcxYaUBwA8O7MJ5w
GedJduBJblelJ7IYXrE/+K0ZdM5aQ2BNUUdoTWpBBDY5j+EGZaGxE3EEbk5O6Wol7wwut8yENek8
xjQEfCtLr6STGFqXTZf3e4woTEv7T1T+yc/sy/irsMe6NiIObmtRgBWdHkApBBFycAaCCKMP8u/S
B6uuT/hFYn81kleEPhpkY250W5CdYdxFBvTOUpD3/+N/isPQ/nnTKeSjzno3hqaywSPGrrxh/Wf8
tc91xFDR/2ShIrE7q2G5/OlEBY/ieZ/xbww4Sjyk6CQDK2XHham+gyOR+aQQHyL5jCoS2NOxw2lx
JJIYdt1u0cUCEqjj5wJOXMfZ2j1o8oUToJ+KxxkSnYQhqRsosE1ZX2R3BwAgYvW1RkFpxGAtdEgI
Rn6/aH6dAnxRhh+yRdcVbd0DfUsLW7n2lb4KXSjwBFU1FDRZYUkSpWBOoH8rxL/F0RW6SZkrLR9+
uQCN5H6DoFfbsA6nmu0ChlIvmcfi1RMXmJ26PsP1FHS4+OwezvsoCL+Yho3gXw5Ok8GPUvCcFofA
SzX+pLa15hQTPPk0mVoDdFug3ABibnxkgBzvjdTshKzl9AJmpAo5dkmicWFk0Vu27iqBNkh3gAgj
sp4GihXX+A//yW/8qEspW/4y4o4awUwKfHuwzmRNX3tXi3DBj2Lo9M97b1zEFF23ozUhog4XZsFb
laR5m0Ii2ayNxOZHQ4iaXKsJuzukJ0LxQYOHgp6LeKKGFXLn9cvjSTXyCsB81kABwBVq4OcLsW+O
P3DktNH0N1rnVjGftXQtvP7cVtsGoIL/MtgHJPSBzKKyNTeKWR5N+RkKYFMlda4+K66DAhTTt41l
3FhKGEp7Bjl3QDDWXgqPrKHHYPiiZseXjAOgFJalOhLWR0t/ce1+nLtbWW077xW7G7/+qNoBC1Pm
g+i7aDtdMq6WR/uztyEWyP3+R6EOAyhyVg78NJNFQnGmGWwn/ouDtyYHhB3OrQBmzcV5Gun1IKzW
3EgmKOBcMBF0gf7bZHz79RFXpV9FPf69pmdIGt5msjx5mMhPfRV5kbxkXl1vD0hpsUXNfWm4j3gR
4UiP23TbRXr6WFOq5uIvbCSCF3enktxTofyu4su9f3UsCXKPwbNzXg11TzB2EnLjyqBlrwR/Q5F6
zSd1XnioG4T6dNqEmjq6cZIgIeonY3qI9u5YcaGQAlng/aLF9Kiu5myGKuSHkxbIbcyYyN2RBh66
RmhRpVqM3PhiSMr95joCqeQ2ebaKG4n2GAdAdxRAafRu9h+4jsfEL/atpf8KwgFOKQ7R5FVpS4Nj
M60frwOirzcgVeItD77PFLSAH6cKyup5GLd+jzqL/rrn4WRGL+N0pfTW5p4z2mZRQ+VQX5D5+NkE
44A3AJHlicXGC2EQEwXovECJqkaP1Jo/7ErFd5PkAkcHqKJMV9STuG8JxsQt1nj8AVK2dYM46nMl
XTwLBMCak4+rRauxB02JHIlwI9YCvL+gIXQAGyxkSBUtK2tY8CgIp4k/2wGGhjo6kX+IfVHIK+z6
EuxqWJvHlZ8gGUrEVTEP46K+S2YPlpyDyWbxXD6oXW6btdoXT9bjLf6B2jK8le+cwgDGJ3St/e5t
jNpoiSnq0OkrKt4RiSTTpCQ2ADeIwYZ3LT/kGSZsdc3EfFgDl3YDAeFQ5u3RKJfT0HRIlcKzhtUF
5O8FBVuuDdeVe5ZqfMPLsZdTpy34sd322jNxyNcqfA5Oz/qAH6LvJ7zUfYf4NEDysaeeATDwndwS
JUs/ygSKJA3I+oFiHZgI2L71IqoKrTmJrzCFLx6KcjhFf+jBLWQri5KaN5gpWwjBrLXBNsoww+oS
keTQcULwXi47CoE4QCboFTECuz++MkjTvYPE890WeFAdCktl6OUCL9/wrvxnIDA9F6Lb748UiJfr
IW1W1SilVYSS+27ilvJVtAa1U/ohp3SmmCtiNh9vVrYSU2XgMJh+T/8L3pear46xgd1O7JocP/tE
DGhOfqYnsHwb75YiFlVTGlLJzm2mZDULHsypbkB2LiIeaDw2Wnxe+s9CdJgBf7VDCBzFR869+yfo
QBL41KbR67QCnHUwDu91jqFfIXwKB+KPIqmSku7/+vejwaqv3J5/t1FhYgGv3Z+zaCFn57WI8NVn
KxLUwUQFzXaIy8tG2Vb7VVt/MKxrNN9GI+xbMAG6bgmx3OvH2/dPe1PCMJtBO0Dx/B+4Ove0EwmI
H0EwSZXt53yAskHaAOC5fvTuCYSHzyVW43qnAAQkD1pN7MRUxxjWkia33sbCEciGgTAKwJS1Bsde
/uwB/M/Tc5hUmTenUFP9nnoP9qwDaVOCXtFXrfqJtr2yRXpsFP809wMGKb1IGd43AFDYiry6Hh8X
jAtLuza0l29qDR8KN5vTsVVkKFFs3VjdxgtcLzKBkGOAlR5/+JqY6vEgMnZqeqfBBQlBZt+YbmNM
yTPkNTVSTq5OctuyGMRpQXaXMl5Io5x+eaEI3uxlCxAApj91dQfT39nXRxs00IT7xwNNratGixeY
Cxm6zme6cwUo7AME6LuUPzWfu6a7ix7jTsaUm0NnW1ZUGd8lNClgk/+9k9MpR80lU2WcMBPqZn73
En8cNVYliTsdyguxhW4axL/eeHjCLww9FKRY3evN+GNSbUmV68gT6yq3m9OECug4mq8ZUqBKTwn8
dDF0eZNlowCXTb8cXt2VVa5IxCi0eHXWAaDITluGaHlVIZc/nABlM14rdlBKvdDbwlSGlPO8BO4x
ci63E41wFxacLoODA+gGrBap6WqORuoPVO163bp7Q9ylwpsJd2SedHQ7Cw/30uA2BLWO1MS+DQPn
BvUW1Nl54GXRGJMEC1fCrXcDSHt7bNrfteiwzoRZJSvhOfcfLCAKOzefGA6Y/JecBlHcZDz5If3k
Kh6HWUQtSZQ++sCmzk1XLJqrJ1gcWLh+5p4kCk4cwvU97IxrtfxPi/rl6Wpfxqpgd7mssIVTnio1
nLtQhU4H+mVOnBWcVhROsC2MegZa/AdcoO9GqX3egoRnQy9ko3+SvYU1y0mz8jVBmaFf3Jw9gBDi
UHWXYF81FIhbC1yhpBNtqUu65SaTd12RB5LcBXNyxHJiXMo5rNjKP8UBeYrOT0LzhFIiq6bT0GBM
IfXlpEYaRGhMrIahoGcXzkz1hG06OlJ4qCXyo9RZklEIDuvnaTPITaQnrhOwQkg9
9zPJ+hYM0w==
`protect end_protected
