`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nvoSdt0LX/oRiT/GlLq83JJev++GCwYPJkLBBjLocCPnK0S2KvlqHr8uL4FmicOvi1zhYlSJlvs/
MsCvjqPnBQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i+rrt5DPWstWIXp/sK2fn8UXcsTY9Sv0eUP7eg2Ehl83WeyF4m7EHHfN204jBakjrCDA5yEjz9rl
1gYaNwgP6PJw/b1aY/ZGWsfMEWTnjxjxb2nbgdFLWYPy80mGIvmqo+Ge7eTTLVKrjMGNucxFC9x1
scUQPfdr7jxehM5k0qg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dPe6rWTXESaStGKU/1pquJcsEQ8+5Dz7X2qNaCEmq6srdxLPSi6P+aaeRcNEU7eK82YkzFvv/v6r
9hVCZxCzCUxdlZ0Q7Zu7kgZCV1qeT0LOZwtdD/rOwYCXpqTYGLmu9z+Cf1QpwrZsEsH+Y85+7obK
PxUcaAAmuF1FNlkNpbxokzOn1qeJckJo4kO8Nb0BQ5KkP1hTi15sdQHGX6TBlWRtY8EQiHZioxIK
FpoviPEcfygIzzSxzBlH7sWhjHAeYaZday8Yp6YU9Lumj+XVG15/5Gk+Xo/uG/UX62IRD8ivfE2C
qkkURbJ/I8TPILn3Af2GuonGoN9PMUACv4qRRQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fVfRPVDBBROC+Gp8uUbD8Y+9upTBtdRtWUOZxTc6f+BN3ut4IEDxWIe6fogeF38DB1L1LmH0rfRQ
cx1fDBiMs6xBBvsgKtgdqqzCds6F7guVI7oB2up4v+ouCsnc0lYm+UCq+QOJAxTqjGoJzrGAn9zs
sIsYYjBy4YPxzLnoH40=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fiTFJstA+pv6KZQynIO5uE4XY92VaF1183uT9IO5lc0Ynj7IfBlHRdRpHFxc0amLoYSom1ceDP2a
6HVisb+IWM8LXwBGDmL1nmf+JvRP4A4xKn6CBjWWcH5j8q4WcjakLcvkQ8HSGlKTc2eT8aKh37E3
kM93lxyXrsCyQLSj6zNKAOU7Jx4XvNcmbllLCdR28ajf2YA3axbhPw4gFYr06TysKVfXDaOZntbZ
wOCIFkstZNM21IAh+JYE3oCgyEYEBM4xKMugo1mkJpzCsItReynz8E+WXWEogoI1EyDgkQ03yrV4
rMKUqQEYgaSMmRyxWSI3/BtSlPoH5WsUuELXMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8800)
`protect data_block
liY2Ngv951wZPmSprKVxMeV2UuvWgj2a1+bxmm8pZNUXYU1bsHrCBYec2aeLykvj5GXLycWHPz0J
9oHubBA5gnsRcrusff2Z+wFV8s+ICtL9hIFj/gb+nwR/h/drw96XoXVMjUPYV75hxfQmsendiapv
sfsdMasgrv1SKj+0KvQnppOtLTZ2CSi2hycb4Ova4IAm2sBn5dP9DnXdiGaLajEpyuEt+3JxZ0sc
OqbG2Fb9vk4WnLKGZzcbSifQXjGHecK65lAuntTNogyG+ggfMiy3Bt2gStqLgmF5yrufntIUegyH
5AUY/EmuDPjuzXmZWSEn0CwN7p7gsS5HXBL90xfLHOGnH73q8jLyRwXLE7MXe6ifgX8jCdKVnvbV
uhis1TeLhkY0vRberI5iMN+eqIVX2EFs/bftagpAoDwRr+9CM2XOydxGKoCeTCJPKRCZkN8G/PRB
xcICbmv1V3p2j0mGNiSMi6FgvIS6d32bZIP9dcugTmcXfB67uBgGTsNE7nXl1r/eGi3wqVAqHlrk
DTrkLBB0E3Ekf+w7aXYBE21no2jqE4i3H6TY3J2hCWbAEDnjeycr/XB2Yk+nRrDHwFkpZ/kr2IIP
oLEThYMjMXdDCzp5kUr82G9RL0vgoCqhCJXoBQIvuidiU5UhpQKICsuZnLXyNzHYdV9DH0tgp8ox
iCVNEI/N5l8FqBIQGqquinar/icbBwSi450z5/wtIgd7ycMJxL9eiwnTxopsx88x3hAS01qjM+6H
d+sMkzenGx6eohneFTpd4w6uZnvnIpj54nT6jCBhsVmSoJXYBvqm1lXpHrD0Qc3ljeRDzWusmQy6
Z4jK26lGeLh09w8KRHX2+XervR/dKnGZYQonpQhAo5Us415DqJMG1dOoXoYiUeh5TvMb70Ud3e/T
qd+y9kh8dFSo4D/aJHR9RbBBai3Tr8ipwYTOLTn8/IREPEZLNZPSkYvORN8jCM8MsRMmKfqjm3Kz
8sQX+4tAUWg6/myY4QvsD/Ayh4V0rHlWN9/yFMxyBH8CYragBch8cPt2KfTjG5eNdvTh9av1Ituh
EZk3acHR2YdGujlTkOyhyXK0kPUELDwmK8QoyhTCdZH9yOQb+31gbuXE2LAQrf0rErTpJvE+I+rs
FMM0lOE8FRyGCwSciAMHUIbN372IzbXvQ5IsdEiziJ/jHWPyGpaydjetZ9JmaxGk8kSEPCug0ilx
LWrEJtxGjgK9p+x7Kz8q1iP+lvLKEe7/6/49gqwjnPjkE1+36fc3fXtHp9wEKRKMTDc42ppyjX9i
g/NSeGrDdtW1ZimRJCieSZIAvZCK6PYfNIMk14JjPmCgbOf+V0/hKZff8Lk0g5VXsVoNaYCh4sfn
HvJKVh1gnQnfPADhEfPd3OwsoYX93jr0jIw5DO86YOYKZ7AgSAXTavZ8NBJvX7hpxQYK00cdLL9I
4aK11vq8ccL4qqGfBbPCI8IfSEdThq0s3KDU3z4DL52HJk/3AUIa3MvRSVwG+QgMk3O1WO9PKamu
CKtbtnfSlV5ucH+TlwnjrdMnMNrcauuCdvTKeGoCb8pOo6y7uuJfJ0e0vdiZr44whQSqkNH1DiKR
/W4jhXN32B/6S/YV1fE1t4cVY7A2LJ4I27XL6fFNmkrkr19wZN+RPhv5Z8g0QHe7evwbfFLX5Gpj
94ujdbZKif5XX1Ym9/ZMivFU+9zIIovgkg5pQ5kn9XBE8ujtDN4UfEIIzvb7gL5vL2YdnqYTXPWS
W8VEhejuyyVW2BlMLoOSyzqerdzJeaUHcohMnaS2/Uj6BTJ09dAnCxcpIdSsUp6wIu4mU5BGoBZv
ZB7sSuE/KQSJsED8MHa+Wg5/eHrFGoTcbQXhVcTImsIQnuLSpcSAHxY+VL2+pLSUuQ/HDIMvnQD3
mFYQ0hymg9OSCloumftF/0624SYjhc02SnASAY5GOmdx7h5q5tTy8LQs0zOjOZuLF1c6GGCF+tLd
tsiJPWOlcHjAcb3Ome+M/Nh/TvVTtN67xsQ/2YhjoxebaS3vYZbWU1FS3CyaZuXKAo/BR8djWA4p
u0mqi0spEEpiNlIbDEFkk1CMKFx4hwe7E2UA0CFXT3Jv6TgP7y1+RYtViOaoLr+a6rA8/kktW9xO
Y6oa9z+XJnK4VU0EAgJrdoq01+WicWj+Bm2as2eCOFWHnz3yvnR/8zpnrbeDnBXvPDBlgNpkzqLG
NxrKSaeVB/eYrLpOlBjSlPgOjbU1GwMOGl026qg6Ea7DN8shEFiwWUWMzCYFeN77twgICA6Nm9Tq
UY3lCpxKdwcaGeg1AxZSeoiXjG4OJDV3kQZupAdox1dbLFRmHHr6uYVzdtY5SkKsqUiJvhYuT3ot
aQrqRqxY6OwoQpOh+Sq+nY7e4WnYZ7Wn8ql2kHJDkAidG5FySphcRZOpmkP3yvF2U6PxdSGIoMT6
9vmBFunSPhYlySEFGFCOP6DXO1eECO0bFN4kB6m/tpvzgVXRxF+EPrrXbNnkkgof1ylYY0uCwKLv
3FqcwBV26wcJshUWqBezjM4nFrNgUcaW/HN3thtU5WdJm0QQ7Ep4Dj9Q84tX8JiZmo+HKk4Q8/AI
ioqqOjebQJlAZllRNoRbFwugtB+G60/Mw4o4DoX3TqKeaoLXyWdvE8EpMzjCqAEr4IoIRJcMzDAG
nDfoNFnkGeR+W/G/pDWQgBuR7VlTqMMbNaH80EF7dsN/FAfM0SvoWI/MVwoTaEn1jxWfK6jrC9fn
ihoa9XZDbM6zXLpnHycD5wfH0JyM1PV0Lp6kjoX8tssXNZmfxnMXPopgx1rd75SqaG9CCGHDhoXr
Invmo2AJPjwR1hYSsZLq6CX32TeOnm1p2SW6eqRZy5voEkTCdEjirKehOre0RT+JPbkt1HqvoEcf
EodrmcczxsjLndHhNdWqlfYg6FskydPj0C9X0AeH8g3QreWIJwR9UR86o7Lm50vcP8RCCptohhzF
TU+JQ30f4h5AK2xynM60RXb+QiecfUpARKEkIRXbAnJQQ9UAQMZtf6AJB07f+oWd9BeMN5Tm/9qy
RPdAL4kyYl74T6m8cHV9L6otIUKAFRgEm0K40wZv1WZRIBYIwNCuQLJuBKo57KW2hUGy24ynB9I6
+cgtvzlD3yeA08/iJv6KN7e1KwMIinfFZO+9fknXOaGtEdBcC3Dc+2vUPIBp4jJtHoF5GTvVof4g
7uud0w68jbsfnHvujQ+nmd78jaagR6MOXb13tqz533TcxFOZrh08JtdyCiH1hW+UnzOKHR4/NG2f
S+trukwsm/sSnffDHGO+yDrOvX6p541VsL79s6USvi75YUePvGo3aIzAg6PsemFlJFB2qXnnWxQT
mW4IgaircY6Tj5SDb6Vp3vUNkEuln4QVOOOkJNC/B/1NEW9AQVmbtQ9vxUiSswPaDWgAevbhje6b
CXR65S19NQeGxwD2hOyOeovIqQNXYpAaCComxGt+o8SINd1buIjX0YM7hm4beTry3gKLNVxsdH3D
IjFxtyc/uFizSjJOeshO9zwJUiNOX2YyjVI0Bdx2r/wjjma+q7cMgJcU2lixN4bbYNwuzqMWgGjI
5TlWAOUOqbpXHpRfXJJ6mSi6eV+qxxQa4T6m0+APGJ/95h3zkIAxB49k5CValKRx8x4EAA8xETJZ
e1lM0rIuQQfysDt2NXHvWORqeOW9AKBPL0x03C5xW4V6azL5tM0wWNo5Faex2E2cK8y2XIlbRILH
7XirmocvNdvlgIPPxiVjpCUb+j4WEKsJdUvG99UhnFuYv5wFqkbBZN6gYkKB7M/aIqx+ysqf1zxC
1Y1/pVVBlpy5pHeYQp0YhZfyJZOP0VDkoGGdbTeZsgpHQ6HxQsXsLl+8toKx20PYuWdFVyfgEAGx
uw16bnx0qSQ0Q6X2Y8DvYCTKKzExk53Xa+3MglsKyGw6671fvQ/xVbyWOfBG8udj8xpj7Rs7eHIl
LTtt9ZIw/oGLZZCBxxXfjlEH42NuQdic3avuQ2Kh2mwJnXBddf+xgc7POi+qAmrpvbwIL7vRx3KU
/mNe/hVkOFHZhg1T+NyrnnMgcxT8TR9Wc1yyMex27xJ3sl6KbJsI2zN6MsNZoqYApxoUL/S9WBaa
cLVSOVDS+BAPlA1rADMIY3003ijIcL2cscB14xO6VrN6fowfb7OZAiWzd/dJBMKttipFxH15fwmA
jRPToL1WtVZ++lT40U4KE/JzaSp3MhSEFd4PLWT8Z1xsSkgvIMDCfON44imzuAri6uJkCBIxHl0E
P3S+8x9zzxWq6T6r0IqF4/7JY8L0GCDfmUH1O6tF4GWvB6DKVyGvVn0xtWSb9sfqSRQnnmaD/KCU
3ovrfRzpZZUeXdEMct/2v5QFL32I2llaxFau1JkeTQzNuk5Q+JqIEMwNO9kLJTK4uB+M+CGhav89
vcypuHkdf9buAWxwGmguGkB5XpQsSvQ4Kjk4BWmUj4dr7cNJyGtlWlow6Pc58BvEt1MbRL6claS3
wbw/LIWAzpSgtQZs5ZsKftMTX/rwUxzAG8yDpOL6WEJ28NNkelkYP+YnzHXzsS5JxDePSPh24gJ3
vqQCRsq0Ih1TzNgwVig9SvjBNaYXVdTQeADrcTVPqF+C4JTXf1G552Bqiettn08+i9U1vdB8RsGb
nj7lqLM3w5qQDeAq0zyXSFmaDYdraALF0/DaVBPNn4QUGdz8B/dfyn5IMsxgt0bV1UfIPlGXF+xs
+Z91M64dp14v4IHClBuRtrk9TgcPliPRzipa8qeRH/rYqd5S1bQjqgW+hR89QjOlZZ2NHyUKPmXT
21AasOiQswocBMbQPigNi18UndT5f0anvVYXXDkGnXe6Rza2jKZJP/cg49y2luhZU15VDXCJclhg
k0VHGH5J4RLkXxg0ETOx4qDfb0GZCQ9Jacpv7OgMbMqnt1ZBe7cBu+2xU9FVeMYq13CE1+CTqzAr
H4joWGuyGIM0aCdG2DcRCd29fn/Yp6px+HLeuyt35DgmI5HpWRBiRXkcCz8r5MWJARGHgWYRu2Hk
ZtEFw1LrrBdrwtGarpgErKY+A6V6+7E5kM4UqBiVWzFalSDnwoyqiNhaJiYmREmkqxG2483lMicd
OvJOu6UibT1P1yaFiFyyB221goBb5kuAPbmsJ2rl2QNybduQB7GgIZn5nwZ5q9yTJP2xMaVHQvRQ
sGqPW2rHUzu4gLsGxF4ORwGMEE68X3+heT8O0fxhMZ29O07pQGwt3LBdpd4iVTK/i5SKXALmepfU
qb1Ljpgl1+oIc+GUS/p2YpdKOkZZqudwqIsOyU3ArrZco1PIhEZly5EFy57CYHw8ZavRRkVDqt2U
wJPa5x6bl6jUyFWFTTiKdoUu/5uExLF6nIGmEkgq5NriQ8fsqe54qRmhPYA3dUZOw5Kw/CUcocn2
CmceT7ZooIGkmXsZo69CVZ0TpbTLwP1zcE8UxvH8r6Ak7AxdWBXUHWuP4ioSEcSdxVrOXOB/08gM
vxhPH3Gs7vDpKojLsvmNdPfa7oXXchi4s3S/YKpiPdQihbmADsJukbCBw/iZTHQGtk8dwMe9kwjN
IB+0vtZSbBG4CSdB1D6o+qoXURnCrZvb9XzJ3H+l5DuYl9yoQ9wBpRmoX7/YGB4WOBJqMKgGZai/
P9tCUpPwkQDnigZD3Jl+liPm3ALs6VF6L9Bd5qAPJ1O/QVvF/4qd6V8SoR52YVHnyntB9WGi2zO7
DLOn6qNErtfDkqnVIDm7q0Scn4mqyMkSkSaPJhy28+iY9eSyLgbGpZkjXpJ2UgDguwoKTYIOqgbH
Og/vHVcMS3gu/uamKXu/Xn9JvC92oMhruuQDKUrySuFANtJMnxv0CRE7EX0Dp9vbtk//Ussj5e+z
61B46GI5KbPtUH+DW8TbLeDVcZ8LGQZg4VXYxCL0/rNx9nHYGbr9hIhLkgoGthZFVrxZCHcg5wNu
bxQllL9ki8tlcEs5Gp2V3qvZQlD39KxOFRrAkFePRceQqzckG+cvSPQED1cyrxk36ptP9b2pcNhC
stRsMMP6Wfzj+j5n7rmbhURvKkjH8qC45t68HO9wp42PfEhLtOJtcoGl4uWDUErDPe0R3QQp6mQS
6bdf6WUQYazuRIefw4N/52dSJsFgIFwPDCaozFvRbK96I91iw46K/DeqgxefdHPt0V4XqqjISLqX
ePNJKtwEHh2x3LmV52BVnhatYisccUG2wL7zApyIOLxvYzqj2/aSEiaRoobhmtd0bRPc15orZM9q
CGoOPYyLqFiTlOr6NojBU2lUJqof/fjivsJyjTyZRdcEXQ90OcbbWOT2M9S4Izr2ZghADjZMu3q3
BHOhgwiFSRzdCcMDouFhl6c+VBgrE8zgBG28OcVMhob3ejZkuEoYkciGhX1uqXSgxMS9CgksO7Rw
VuU0zT/RwuLqsa3TLqMXYsR3i2uT1BmEkUXmg0mgF+e+Rkzj9LlBYp+Uhgy9Qx8dYqarcQ71pgus
os1C8i4FzKwY1Tk1N7DRnWhMbBWSB+ABlUfbDO5CGmMDqArhh9vzm/QsYZGj023IFSxslpPK3niZ
whZPGQdyt/y9SKuZwCb7JyZieaK9ScjBiaLVRkZQscrD82809pbms0XRW9cmnMght4Yf3waFzm6p
M3xuNJhFm2vWM1doJvz1pTlj/St9ugQUwQpLUim3NBGXGMfetsmJgYnVIwClR6/cTcCJ8K0hhkl3
4ZOF+IOwaX0xqKD0p2XbK/G6Z50c6bDWtCNVtF8Zf8bwiKQ8R33X7ENYjp4NIYBdIOXvtQdlIwtN
4UqRM/bTza0neEPl3eqNfVBOElJdB6W7/PjzJpSQF/hNZhvDEz3i2IZUEndVy7RideZ3nWR8BLeW
lVQGow3t1Qg0i86ocrn4GXQoO5nbtZ1Q6HsSPkmyK0xL69jsHCyWZm3hgLTGpsYe4Ma+oh4SYsfd
APQK21jlp+MQKqRUR9npjgHe/FXRrQ5X2GDb6wpVJuk6CuMwStunbPS8lPQm3LkCPc51cPuAq7OJ
nC+a9HXGpA4kt7dX0moxE/OzvGPwJte3V+Q4gReY1I9dllm7CApiUkS3ZK/xMMRFAXHCCSFWJaxU
DaB3AINekv2bIA6hGI6U1xm8TII5yWW6mcTcCOoqDo4tfELtycHZ6yqUOMmO92giLRADj2IsKzJa
teFt7aSZjjgT/AQ84s0DOAKbP9+3gTqEwEc+wt72EsXJqLjH8Ww0UfoORFv83gqpAJuxVNBreLii
3h5t/ZN+KPKcPOfQekNoyVXoPoUWIVawzPofep2hkJ1zVjvZ4rTwXTnssgFTKxOr9tROuDF/rY8/
ps9CNlvoMykG1iC3HzJ0Dtf7jfsEuFyscHB2kloveqIRfUCiB3dpXfK8JfL/9eHqWq9hdvWRraKH
fJl3hTg1Wsk0Bcutvf5Urk6GErBSEXPGDEkxP9Yz2a9SGXTyKXCkicFrerR/ACKB9JTpr19y3GmU
ESTUib/CGv3EB18cQ3PEhC5GCHe5vLG+mNX4smab7xphIUPc8HAx6WN/8m6TDNq4udxpoISoPpYz
pkn34flyk2AxC+cKueUeL8LlbrZoxF8/ycSLa8cKPJjK0x1+0Hg3vjg4AE3sk3kAMq8G381cE7Mu
V61/KVLxyQxb+3BdZUA/rGyF33xZxjnwTGBWeOENWcACFkQZF9+JhH1rv8HmyIGxUhfYRYm6MT4l
QRPtkl9l77Q64ifUxYRl23AOJsSvS6+lsiD96gvYH58CZPm8NcAr3nv1z33gGvVuw5P7cX7WcD1L
ppTFTTLtauHRMaKyYbPBqrV6TrqwIfdx/wQTka1oirmBla6T9zG42SBI59jm9txaIUEYKdsobyNd
zZr0/0Cj7V5fe5z0eWzIc315JMXb0cu4P/t2+V/6kA8ahP88U7kEpRDa7yX+d9pbanuSYNMUdyM7
ax/sDS1bS3GocysXH9xU0XXK81TKxv2C+KZBd8T2u1X0jxoNMx0PnJ8omYiY264MTgfKh9/t5SU/
s+x1+t9nOReSpAzgyFFexwiiQR9XPIvPy43D1Ifp3VZwli7q3+fJbpTclH4icBf+hlpZjK2/L/0L
YPYWGQhQ+ANIAIuVa7MMqV9Np68rfp550E6zr2w3QmEUria9zrPEdJ6FhQ82GqGBWLZKUbFr2OXM
XEErpsNWSSISTNq8yWuVnKCOF9XmtFeGonrIyh77e3kg+KvwtcSDzbtM0OVxcM33ZHpbf/e7MEkf
1VW17EX3qQ3zJK54IWG8x7sDijffP/p2MzZ0nVrJn3G19XEKn0drC+jvkRsHTQgM2wFqwrDLMsbM
QKWrNixVb+iqqcLfgI5L+s9Go7acsRUMzDW7GnpqDVZQgj1n2szRZk2IzmlSveAQv6/AeVgE1mFf
cQm4b/eaDWwarFViW5mD0emoSH9+MxTJlbSUwHP/kwJ7cDaemodrQDU47CV8dNlADrlxfNmrmeGn
I1osmsApBAuhXSVaei80Mf6QwzuyNtJRCp8xdq4+FccTOEPChy95XOeh9EKqFe7RuJiTyQoJ4/kk
PfqpvZcycsLOEeiDA9XbUGUzn3itJEEzFZf3D8Hu/wlCToJJ4rVlQxG//1YODxqcDM/v9RG0auxP
X7XdIbpl3TspaRr8CdsTOmKYZC+IYyUHwAucciRs8F74x6aGE3dBFCmpGMFomfAnU6PoYZW4vBuN
/dSlJCaCUDXAIGWg9D9gW4sy/WE2YG5bWCjXGruFlAKY1YQ94DkRii3MD1IEHRAOyFWhxnCWRSCx
YpRb5d2s9M/b84K3RngOsQeqx7YrskYjvAxnfO7m0n6Q7viwb33EWOXbyLLEyvLlHp/WzBERtNZK
jcZpBTkBgcwihCUj0vQZEpGcAqanQ4Tv807fwGy/QdxKz+XAo8cOtoeIJ+8sKp9oV9z9H+RmhH6A
YcBQ00TfEyKwHoQr7a98st+78wtTBBHrHeefwNqyjcb+BevCWrGCaKtTkqbZ+xoQy53Cx2g4P7ES
qMTdJUbaqvAqL7FWyKH4CfJIodR/onx6sy8XHqd3V4DJR0Zw18CFPp6XR0SHIIvW61XbMcXFWKU4
+9cmSHoU/HHpfeXbOrvz/qqVwDjxL38L16Z5aUgxW7B48ZONuSdc+Y2t3ImrKmwXMpo3fcyw4ofE
ku5WxSFw8pz960hRcEq2AyNJroBG22yaVhA01HDB43vsBGwNnDqbbhFZqur5uM2ycPSXTo+aPrFo
Pef2Pf0QIq8o0OatrnMvdp4W+t3ACOzMdeC/3HdrfeZtCTWD17F7rWLwXdlYEpLMkC3m5SOo6wwZ
hM2LgMJ/NkSdshO0bybYlkwUEGhU8UWpgiGTxIENS7GBOt4scSKXmc81J15vPeq1I8gRROgbh4tB
mOmxY2kvZ/L2zx6yN1kheYtSEudj39m93bWQTBjqqcN/rE0crkl7j0G5kw8NXpDD0RYfkGW7eKtd
swlslTj3sTdh+rjsnGNPrumNgvqMLMTzMnQv2AJcLdJyBRC79gXM4HtIDPkpYFS6T5SIgZJSxWXP
GzUYkViC73Ooej5Mdr+uFah5kZ/EgsvS/Sbr29ugV2MPJ4httpsZgNghHAK9wYjghnnZmTErJ6s9
rMWbEc+gL02bnHAkFpshegtG6kshhTdbmKOcWcHsl5JNutw3hYpZbo7no6ibZN0jD7yMC42Zh5iB
YIfBYLpebA9UQw7OFgZgg89nmggF5dpJyrKcSRH/MKEh59YUsNgVgdMka8/pDsdROYomG1OB005r
+6dkAgJXzGSONsqcH3WMqDU+75s+UGEjZOSc+VEsAdD9fmVSRcHtPohSJCP5dS83Zz5/AjHdS541
OuMJAFbomTA+tfr4OXRjCHWZKTi4CvsUyLu7COhT9Pop9/n3cWMz0Vz23zuH8CZOsBXl5hujiphm
b8KFSzVOPSfQXk6PvVFreE3PII+91QItkTnAk8EtXsMSZb0yWFzuZ2Wmk12o3sNGCsehGb+lNTel
oU4f816w/vc4iu5H1Bna5+BOhQVW65WGaXZ0cchyJ22ENn8AVr7FQn2Hg+9OExqo7FPKvyr7zUpX
clfR7SQQBC0ygJzfZKhoCvNn5/LVqWPPpSUGmP2+kD+KqJRwr8DANeeS96wxQ6xBHCXRlAgvOTun
RhBf2yaq63cFi1X7Z8LHMg+DoTV/Zdmlf1sZnw1q7YCRNsR/7j9ItYmHkIh/B1KiAu+u45u3oKyg
XskYu48pNvST//EOnMLsnw2zSK+Eb/voFh1c2Q5vGCVFbx7UdVnCo1MHSp/mZfNI+Nb+/dG7kTx8
LqXU+UULnnLiHEmgHbRYdjE+RSNkD0jdHfzTb1f+PgN6Q+NY/tyi/q8cSoh5t61KEJcakETDKObx
2DDxy7DUXfF2S092KZp8LVCEDKpxAto+WG9FQgAw1kqfgVfS5GuMnCbeKXFZIZFvnNkkMCNSpQV0
pWK6Q6byh6iTxI/s4/2TokersSICKVBT37Ipz39Y3A1We2g41YR0KFCmYtTwCGEjGCZZbYGu9fzt
G4nMcXgBOV+bAreD5yOY/NjZInmwKoYCQDMvkemYM8V6Io8B6rhTZUaDEPQ3OdKvj6GiINomY1u2
Z1hsfB3YGeW4FT1WU2ztJO5WGOHUVyL5ZfKg5VI2glAkenkj8sme+WStR+vuJnbJ3iMSDLt+119O
wOIkIAacfFK7N9TsPhAmJotnkzfmUBBZOSzShUZ21RT6pXTPjzHuuyCKViJJ+4RW7vRHyvnB/qCt
nRO0mdMshPGh42W1oVx4NI88rDocX8teGwu5TBf7T+3fe8tLv01FC+5YSWEANzSMawxSW7mVJW6r
mW0+kdb/uudDt6bWSI7LVQCycyYpXPrDrqPOcqqSRnZ5jhtiS4blezAnUBMw+JW50a70j6iLhaEn
xb9zkf1UUHaR9q09Tm3Cy4OqVF4EldwZOXKATWDjapZh/ygiXC2GzA69BmgYQVHbuDyrXcZc3xTb
yvj3k9rRh04XkdOP0kZGl4zOImPA8MgWIGAvFenRDZPOKQi9456sYevjAgjIQ65Hx5vJFBeH1VyH
MxT799H1ZYuE9Y8Lh9yNp9Se4ChnhwW0t8pOwJhGJF42AcfBUxRvqK5+Qb62cX6iisQTJsoPvd+Q
oAFSVXCxgfShJ6AH87IO8gW7MLjhio6bFukJ2q+FnXYL7kMZ/m5dwsD7S3Mu0s5fusOttOmg8u5j
u5vPJlwFYA2NFcccmgM2z1Vi6+x+rE1ghZuD4QPgcyLMy0YOM+wy0WpPBf8ij3CDzNCNbw9xpeaf
P+5V3lpeNkZ8EkMrnao3yHFhrovWm9Mk0aP99OhBayins/19dXIc9Gb88fhoF10pA7OVoy6NwtZJ
N/RJR2tRcXAAbtwkbByJDjo4Q6xAgNlx/77sJBLpZQkhtiVMuTrWFL6IFaFZrz+d//2rNsIlBFth
WldXC1t2Xnefd3gXli+xCSORb6kfSRYR2owdxgU6t3fsS3CEOL0i55zaytZnKWrwaZiwqHi5pQfx
D3iNiwwUEmeyUsPUG9xi0gYBP6rEYY9yjFnxlv+4zD0qtGQFy13AK+dOEpaqIqnQ2p0401zTsivH
8Nmsxvs1rXeuwH+OegkiudZAuzqnXF6kCq/5z6Y5MgGpgwnDD4xPl4E+R0dCTHd2o3It7p8WjIHF
fubijhtj7YtJhJelD+NlFoMP7K/ZKjeQsDMu/+4CgDW62uLOSAr+c0Y6Q/l+zLxxnGXpLKu6q5jK
K+XzwNlcZ1dNjAZkpsofmZ//vlHaQw==
`protect end_protected
