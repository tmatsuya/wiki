`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HacNaRwZ8KPWtJeWFUwq9f9dGtR7D2vf1SN9S6Ciq45DgXPAlBVgHTDN7v74C8BvW351s6b6ovIB
qsujlvYpEQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NbGYL5XlNS8a+2D7yDhM0b47ke8IjHplRYKFR08LJMuKKqa0KSBc415Sj60YEJOv2GZPIV5Vl50z
BphnkHeN1oAdKLhQC2vYbLUH3DjBOoBitG/JAAIJrIdrM/ftFjwin6lLPEtNpTn0MVjFdPCfrPS5
nDWvcNoQuKgYK46urZY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KTEc8osKqcoinX0fUjAPIjfykXMXU0j1ENhDAccUcK/x/VSjp3a4DcQqY864tWIhGl89sVkTWtgF
FpxmK8VqHWq5boEZSxrgEN1aCsdHqBdELMvwayZ6HRzjILvfvsNjgoLqkV7ciklyKN36hiFXOkCx
WP7ncX/93RGp/+J/mRKcSNAVQf2jG5A9YX5g0u7qkfbCG3BNY9u+jHFzerOqTDOjOyEftePeDEPk
7v9F7JtT1twNV6BMTKEB6yHhnkfwmu4kBtHsXgHS0fyJDI86x3hRtNTSAGCghPBMddo1oUzbqhia
4uGLjzY0XGvKqvpQULAhaDChRpNFDLcnJ3/GbA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YcYfdVgpd4qLtZlODmK/MvQah+Wf/KcLyg4bCT362d47vRGdJ9F0qvCr44nAA5pIMB0trrzhJIZH
8a9EFMwrAMfr1Nkb2RVM6WA5IpVEhlSkTPkCcs1YUwXH42DsqAparwSJS2U3nBuXDTM1Zl61pAGT
0t1OlbKxwT4vzDMS0S8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XMXqvDgdl0sgsmD1QfKYF17wEsvKuHC3jGY49jIY42AhcH6H6KovGdTxfLS3C4gkjc5XUwXBml9y
EWllSQG8GBt7PkXO1B6sQu1MGoq5/7esmqeZtrwsykcxlF3NMT56kvzZDh+yUKGzJesRPs+ukcMG
QH4Om4HBRlfGIlfbqlbzjyHdofETKzwlNVf97D9ArY3yXbupNtU/Vo4xvKyX6SF7m5aoMxCR2I3f
5r2HZo4ONRJ1Y4f0ZWMDHjTSrJQ+SaeXhC26GHAIstrbxDw7s3x9dihM/h8sZaddurRBHSyyBErF
nlYXqDPv4PvRhZYCSjD5UvY6tZs0z5hmQ90Oig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14976)
`protect data_block
xEObOWA1dsat1ZXG8xVmTwkaN/yMWXP9LTlSEsU89YE/Sx9vu1RAscHVVUHDdztFjp7gweZQjAV0
IHyOUxVMZE80NLcdPl1jkr6ELukJPH/GRGa44yTjRoyZYBbrG6lcwDvABkl8jbwrV6IydHnZGG5B
e+UOly6iMiYMUx6a3JvF1WlcDhAchJEdCmyuvPOQey0TsrKvSDTthq7bJgRRIrH/A6CHiVKMsY8t
qRL1UsR3jH7W/2xv4u5Llw/ePpVkIlHqGIYVYOAeR6x0ah2SfMApt32tFwu1+tUDLERYY3ThLvZw
VA3mc++KT5uf7SlrfIKy9Yl2MaUT815uexI+1pyKaL7O1OnlOoBihacSjgebCT+N6BrNDPx3yjRx
p1yHHxQW7Yl2yt0NuoU9mjYz00yz9qxRJt6Zv9GhkBhu6CS/qDqSyBk5kX7UAn2OXJw0068Pyirj
BSWDWU2z+3FRu4HSR5mSW5ZWISJ1lG+KJORvQite4QUIaJBMyVYXnW2Nv/HXtQXjeGPTeT9DSZ87
cnNLtiGFgia1w110hH7kX91s8MZNJpGgl2wKQwK46RzMKc61n2MN5Ul1rysiy4gIPBQ1cm1oxq71
gdW5Q1GKNS0SAutYSTdkT2SMMauu6G/9gINr01ngOFZ2SGioUpMBH2RFe1RHNUz5WkD1R2Z5Z8nZ
5jDGXnPu+ORGfSZl87lstCG/UYNf8RlNvk7VMFTq//hgidtfn5g4MgK4tRl/6F3z5vo1y0w6NFF0
GKGTZapRupfcDt30TJNKKZTh/9OFdvUe0rWuxEV+Nl/BtLXHhjAThuVAxo1asAFQmko1RavmaJ5t
FOqTe4PHH0XaEc7D7TphBlMoMwIOkXjfBZGCabtTDY7u+EfcYp2o432A//LIE21Sah712bbShs1h
84JGrqyYHmbRCdomDSoxocgaW18D4vNNNcKScUoOGikmhXu5Klg6nyTpf8Lugq2DU3A7a4Z9CJx5
49Nx8Sotv3iDSqQAiGaJasaj3av+yJL+0GMNZYjyQfTZmSwIhldAUDpd1j3VB0dZ//iUlwSMKqcV
My81S7w5U4AewdIupV1y216J67waWbXrvoueA0V8w8oYdUJpCw3+pbLel4x+G35HzWkywXp40/Ea
OfJDFZVDdMbpudlYoJG8h4tMv+KA6wAcbhv0MNPzCWgrX4TVWmrrWWRr64dn82PIngNPdlfnbOzH
6MB2R10rM4gWRGm0X3A2DCvC6K2VtbbrOm1W+41cnBBwfTOD0FNI8v0X1mLoRDefvLpY+RiToKCb
UvDMRgACIDp7jFTLWbyrm/OJ4ppMhvDCVYumTUiOMJ78nSQHFdjoswljRbgk4O/03XV7Et53u4pY
NddSKTdU33T4fRoOJTlRIUdELvtVgg6uOSUtm249MlKLc8h0T5Uf8ZFYuN6KZ17R+Rz/FPh0QdAl
3xK044lxcg6BMn6m9ByBACGY3cKkFTE5YhISVA1osYgnXRdeiVVhKZkrTwPPSNWnwoG8YqhdtEdA
KdWLVNhN84ATY2UaxwJRf7TarVVV8pBhhC/C8J7rzgVmn2c9fSSo3hftKNxiB5blRCE0j3GaAbnU
/CeR2sEF65j0upzurJNceJl4XbhupByzU1dOwgVl5qdSSRhFHJQFNCocUB8aLPerb7KacYuGfDDR
uTnB7dyfR6vfLJKXKCqRBU8QrPIjzV4GtX3s6Wga36CF0GFrL4fXQxSXdX7I2bOGvmg/aPHYZSjL
sjvQC/uuUwHblWr/usaEp+wKpyZoMh9ZWtr+FE2pjtE84BUmCDzLnG5Ur23MJ4l07f7FTOP0pgjQ
JZHyyWxtaOjbiRjHrrbD2jQXEU4XZkNYm9qiVaf5P3lS95jwTD0uWIxXcTP2EpCzDaG0ZqfTslgq
Ku0wYNvhrHg/dXyK/LWOAqlowj2J+HTZDMOp1wxNRzIHG1naCRDM8idjaAwyJAhfDnnoFBnZJZBL
tsZ3gz6KK3Zd9QtU3kijTS5UCw+A1vOqan0w4zgvcANqD6xMskcLFYJu18Sd+EjcD1aABE0ZshrN
fHj5sK02udKY1GRX+CzdWtyg0OglHn/QVhM/oQVyaa639KoxN6c2RLCFe4OGLph/TIq1jnke7iDc
BZy9pu2jzCnstL4g49ULvo1Ssif5u631ORIBQtOVlsZqKmd1sRTNvr3SwJFWlwh3XCkcZq5H+SZM
m65SyXpzQ9HF/Tdu7AhaYWAy57UBFoRB4uVF5AZ/mNCeuF3u5cMaDgnDmGoZ7bUQBx+aqc5Mqp4R
B6qgH/dOTf8xKq+cJToewCsqyGSNpx7dY1ZZClyWBy4hrqHjowlnk6jqcTLsCzpNbsEGzE37lhkX
3YTwc3TxXKUcN21TQq445vccqrSWLIBPOTSKS5LEpY2oCQ6uKftaD/nCLtdpKfPvUu5fHMNeHryI
H9s1sicuQOL9N2pups71kBupfY2i8FABnl7tC3pGS/HCD6NoaQN2dPBwy2zKByiyZ+lvMVfMVrL5
hAUfos9bzQN5AqysHFku8UhaSlvuEMuXQAY8e8FbUMR7WUSnyx6ERCy+BBMzNob5DkSfnSZPSSMq
YQzUr0FmHy4DbpXEiW9gdhlpRryI4zp6XtodLAXmRcO8oGpZnaXYUvU4I23uezt8O7oal569jxGh
CX1vheWruFUf9ZfZ4jBPlytKq4coRgHsoiiZS1ZqfLFUfC2nwyRoDvEH3Tc1FjtNc2yJ5sKimgkQ
9gQYvV+kW6rPF1Gfe4WpQsuDT11CjWNGbhsMNjGGJV+w09R1Gjz2vBDispdpjggZk7JI+dPYUVPG
QRkEzQ/V289l4fDRGKej9LkI4zlvYGQR9WmtQnnTpHIsDKp6NbySEtAdS4rfE25Hpe4Y2s+RP5hF
ExZURzo1Jie2Gedx+hJq89gR+OpQ3zT6bPWwCfEA5BfA9TUE0XY72Uppy3WSsoOmXoR/Ealnqblj
DkMAiqZg/B4cDyN74s6mWVUDe1GnXEZpIKe+dPiWN1cxowjt1BaEchZaIfZ/0kYutcKj2CvB2Q+I
r+2zxVVB/yMQo2V1e2zmGSsi7K5M+pIa/3x9U7rv4xheEJ5AlN4z8Zmw/4bVjoC+nxmD5bM7TbMv
2z8TF0ENA5gz5uihE/g57r075Hz1Ef2oCPjg1ni3K7FCa7tLzXyG/ewmZlHenU7I9RXsjf+YQw4z
/AlqZoSovta1PB6jlIW1A+9OiPAaJzK43mqq6zoX0BWMSwp7FdNO3ag8QbSAeuxj3EngZ3z2wdBg
bs6Aj5rSRGvuXUEuMPCNn46PnxSKMYKgqXgOCM5v5t7UXyLpltwT/P8w12RzlljxuHnzpVWk+m85
/nFPO0wsFvskXhqTzmt2ZKRYx8n3rw/dipgNuoHuF0lYCjr+iDZfhPOrS4ApgE+XEIKSvgy7vJgw
srAW1SxNpLRhWVEz3yEFPOiyCmuqxJQvCofEH9Nc4OhvPf3FVsE0sSmM3xrvd/LXuibnCajfU08W
zMGtBYoNQ0xtmPfVEqIlKZWMxwHVB5RzWDmPA8esFS6ta5+igiyjz4u+PF3TZq43ThZPYY7CrlcZ
mftMINWtubR9VX/QkAgDvtLB3olYZ6j6ShE1aW7Z9zowRsek2dJAXGM6TJdblRflcfY27O1DUqUy
xhu6/pyi8NlrpcXw9hZr+JdSxN0Xp3ACiLjQIcqZDnw2qeRcyIIfa/T3Ppa71siFsmwmY1Nwe1ji
Rkn7BwcBrR3btvQZpoKQRzqtyseK06kA/bjDePGTAuQ/rW/9/Nnm8HIgLmgd02Hx94xd3OPWWPWx
PD27jNajN4u3ImbOZcExkoP8Yw1F5kOfMgZ7aMLhPdsrf2ihY2cuM+y1E1nE+g1PtzzQ0R2qbsl8
jsoK7vrnLJKe9wKJDsUWJE9UMNZaOrRGdIWTPVHSqotpKCT1crB6dRQMNbusCKr0KL1V8Yh2laJi
VNFWwnLq2NCtN0O6vdaLYUZX3upbk4JA1KqxOk5MKuoKwPyGEaFK7g9OCqgYm6tKmLblNtmjSjcP
MWJ7m67m0GIuRy67mwTvnWNwAE0gsz2eslnRvOPUG3tje+bDEH2ZbendXDZmCyJDGg2hb7CAY1yP
WWoFL4rLe+Wj8oJSBYPA70512WyScdDVnxshKssrJ/rQgQZQWOlnTKN9N4WFqxsLM6gJAZrwHTqS
/24riP3Pgse71I+KqoMPVc5tmMNDO2R69Nj/raupdJjsObMnNrO1g5rcsKouHIELMm2Dzzyy95Yp
KsekraBVFrkkUo4KeBIM/R65sE7m137IFNrMEfbA7Nz0S5h3/OSF2R3svpdZBqfdzEo8HUb+RNzK
j2ICYQo2u7URm7h0qAqs0cg3dIONz8odGw95qiBCWmUcI4sGekkQ0QnJX+Ej4SRYXM27e93b/DST
jKbszvbw87xRNeLKwMHrGYBn2pGRPeZ9GLJoBL3fQ73dSkI+8BM5kKE1DOkSW1l3t9pLGK4DtmrJ
KwKu+NkaRLZH+ICtU8wAHQqNJomnJDxMjiC5bXvrJgoeR7FgQePEerMKiL87myCBlR34KY7WSRL2
I/uoy2D12z0E3lcpsxzAoOBBfk+9oFntUplgaVuz6V/KqvoU/r+znDNHTl1ayQ1MUOB5Xxw0oRNB
Qdg0ZyuhEj2zuCMfvuWOkGu7bTyRQf9xnMQJiyv/0ug6g9D+XtbpNalmcDDbvG7fwFKp6VreTk0P
z6jk2P1fQOF2kfVi8yetRLoSN8I4L+SXjGea0UmxPuocDVpO27/YInr9VGuTVtFP0cAjGm83R4ex
oYJMh60xqfsuGGz+y8DL4fChqyXOCOk8FGwWuHjlIAekaDGVHIevpWJQvtBlCjT99S5mBcatK8qC
0ftzQt2rF47PUaaojoJt8fl07WCwYAjMquJENhQu+XUUr1b1TbC1lPkYgfljJCpq5jS72/hNgBiO
kFDxEtzIn7DZ9J3fd5vwLFyArtQv0TBFyYVD7QLIKGlzJnl3eJK+htsZosyTLnRrBcwskSVDpSmN
08ANYm8KFKakom7qftMIv5q7lWyKEURWeFbNOMGoHkK9/UwKxvCQ3A8UGUdALJaIn7glZPKTu1Nb
kfkVgEhOQecKCRCHpGoOgtJgy7q+UxUjCH7YmVNlqzXJlMmM8Cxs3mFzSWmx2lIVRNzBaKWOxZS6
3bcuq1fs3mV8SXCkIGJIs/Srq0OL2cpv5vSdtNdIH2fI3dogbzLLr1aKoT2FKuHldmaEdxjBBQuq
HRW0S9xoSiSGhKi+6BR8K/wGwXZuWHz919Eyxa5vCR4HMzXwDtgBYCvy61Y0iNjH0dbr25MxpcDH
9MC7g4JNX2tQd734ZXEJtkj8OhbHOT2kZkT4C4JpqXKMCvJjZ88ovxVXgx4OHdA843YiI5pNwjzd
YvntfKd+/Cr6igrf4gPsoz+rLwHerfFk+OgmzFaztiGMPwI1+qQr1WTEXiNPgOPiXjMdgg+PO0N2
Lf3CA7WNtR675tm6TPLGoDUWRQZb0lSw8roCaehnZ/K5tquzFmSw2rgW1uiWgpwYASDp4ylxrchp
HC4IsLV7vrgfan/xYQJRrXP3IqLLMjROgE946DIXFH8cIu5pjVJUtX4Vky9LP7pGWoecuwYkO2tK
GHGSgplZ7mLxsFkRAN0mpECMGF1omSrbmy8aGveQgfY3zbbnbOPGGoP3QW5km1vUFOCWstHI/WTN
zVKjauqB6ppVpB1QpqUKKj1JtrEdu2Adp3eNwudjhiwoldD2s2fj36IVRRht5l+PTn6FqqHSQhCg
v0b6mCpKpUp6G17DwtMhJMJP6nMLrcEt2xDhF+MerxCGCTDI4+s88tGsW4XhJqWH1Kbw8YH99gjQ
vCBJxoLrz+9ZVAtaGXUxoXmMjOqSXLiWt+7Gz8AlI55oVo3AMPl9OIZtj513eTTVVEC09Od9Cxcp
Knn7gEuAvjh/jtHsaW41t4AblWCNS/Ren9bqDyzCv3J3PIE4v9EKRGiK/nfYeT1Fpyg8+3i9nFAH
3HcChTx8XzI5LN4wSemu5lNOZBpjtDVk9AHhEnFJ5gUpAiKYK9dTLtSt4e9xYnzllDuE2DhpLiYQ
oCgd/cf7RlH0pAsIFHpRfcUuhuuhDwWWjLvvv4EUvOxtrPWUZhN/KlPYK5Z65/5qMZMer+nIEvnC
+Or0ZFo++tP0RP4ckcE8Bxez36FHXb2vCi29hkeEc4HHDF0HGTpnaEO8X6imKWXEtgVvUK0JNBHG
R1JR7TYMWlnn/LAyOH3JpbqWq5SOalXfm8uoasA3+S/8U+5pvZ2usMN8yGw4BU9RnUVLB+rIws3Y
TLYehc9xbnWD/+jfSnK+a0VV+uTkA4g+90lHRKGYDxqqlD12VjvSl0kKYnKr67B2Hp8zrLL+OZOz
gSMsYXuHLGNKRsRn8r9dt3H3kfUI8pTUesPfxSmIfCON+Js84I890IefEtvJGp0WEanP8ic9eZGM
yVdouIxeSUJyex6tinTViH5EPzuFWoQ7oiYN3HzsnuocGxxjidyoPqii9C8i18nh3WBNH/77zBq6
PyLXAPnaSueJb4Ach2szOVlpPo3dW1G8oz6Inw8dDZXWhOOqKw/E5OLk6zm2h4gRlLN8cV9PH/I6
dOKOsIYBu/YYEs+0rhi35nWQa1+yHQAUuOyicrD8hAYfAk9ygnlPGyrC42EDGnxUCo6izeb2R+Rf
F2bP/Snpj6aXiYVR3+UaTPkkT3VjYEX/mKucKS2suaRoqTbHSHefY1jXGzA88Faz01DHX31b5KE0
3iql0i1z+2Ccs7N8ffBQgN0RAE5gk2qyReDc4gWo+QHSWXYhU24hhJcOhoMcE74h+lX+e3L9dcR/
r+snYMLsrfm1W/4+tiIFPPxFhhkTEMGIXAWZGaoY/mwOv6aiUSY5l8lgCZ7ZeVxA1ZGx9zxW7+Og
qTjyqT+gMh1mJ4WnNnN9TJ5lk5lKWEexxs9yq6gD9aZ3vMpwPG2t6+7ymfHamQ6AZ8qfeRz+aZrN
TolhmQO23mLnnBm/J77EqWxgbEA7nQbg2xztLllb+lS1asg8EBR0foxD3Ppnr/pwqbWFTO1KrJXT
TGsSwBHM0qZYf8204o+/FHnIhE56njmNVX41qvYFJ81CeA1xfGhVcKrRJjK98+nfYA/U8mygw9YD
ddg35cxvnQR8vLm/UO1vasAE15QmLF7n+150G5DF1b3P93OTbg3QuJXVv9g6gGcyd1cuuB24kQFz
+v1c8q8UtURH35hJ/rjQ3ube6I7QovNNC8ZaMf+v9a1ir6T78qONTC8kiNEqclD2YJRCfTKsZxdk
bqgJGlWQVTJUq796C7bVs+dmVpS+OwAeBsfsNZ2XHJP/kPhxY1ZdXIx5KQBSUcvB77v7rXMToTMl
j3iJueEnZXCc66gO/9Rn5niQ0WQrU/7IPWVxsg83Z089+nplbiXaaK+VScw/IvkBsV9iPjhBqrwW
YzzCHCy0oU09ly73Jfb27Wk3eFwLw1ELHjjfT3hV6r/eH//w9li+fZv8+pOOfEyDhgJYpL+ZpNaa
Zt4s1nqyKsmuCF4llZQPpSZ1qsMMJ26Fp3U2arG1KybVc+vW3oXc0OD+YEDl1rWP/ss60Nz+i0sy
1wqATLWWoPqDcD3qTZntdfbVuS9JJt8ygKf1fb/ns8gbRVdmVDcYjQbkDojRoUUY/C084coYvZ9o
bMnYk8rrIHIGviXvm/kkgj6VFZVGuvCySkyrwEMP8DXfZQ3UuLwdWPXLa1g9rxtqHKPxKVpoaVvX
nUzquIb+lx/coXJNm4m5GB8ZVlcx2344B/coMAhxsyixkQZC5CCInQ0OfysarvGtJyNmgS5mRrFQ
nXalJFHnsUNO5fp/t8z2/Xmvw2HPu0ZOYaj9WKdBoW6C6fR3nk67gm3VSdnK+FGxTniBN5/aqE/J
5bo2G+KaPoLzrXlOIL8BVww4nMuQVkXnIxt+RiAUu9RLCfr4iMfCbmKiYunvpTC70TQnFRzflhwW
vUfDwdQcr0+YjV91R4oIl6fa/NGZq15Za1IzVA0ewiBuqyrRmdmlgZacB8O9hauqvzUhtF6uVwU1
3CHyRAKQHKCnUTpnWPLHSkV0CRyE8Eg9skgO4axMJ1qUGI6hMWxXBkC4wYEppySaM0o4ebgsJ22v
z6SNyU+dGzIsSIjUjEJQDXE7LmYwEzCI7Cc3ptXihUmLmx+i8ahcOItL4TfM2odUuAeUfn0uUZka
sIdq+cwminh9lPo9aEYsXKtxSEm8o5zagLHEqPF5fFY8kgJsWUVIHvEmAiPTy7SFlxyXW3ixG6r9
W2QlLUrLXoIU0XmhorlH+OzAEIjWyUAbi7SscdPJMYRlZmhMzP8dJRKnDyl5zu+M+FKQVXDhxShT
SjduaryNyGq6HvtVI7M0syGTLY+uh9ua4g6YlEhFm+xSa/2HMlXXkunmnexHUzCOAxICzdWK8vr+
6OiXkwZ0E3QAh8lLzpJ2/rKCgBrI+rWJYW6lkWbzkrfhso0OYqHzAttN1sbIGNeUnlHjKuOYp7gP
RSAs0MwcDx7IkNJfZIMbviv9ByUWTnXyhu1HmSXKkSKnmjuzU8ivV8cOICatzUSpt0sQhxI/Ruli
rwqzpQRwzb4u7pAt4rannIqUxJjFiHuI060VJEHLC7ys6bS4X2SDPpjRvr4Zt8MEqpEz/byVlxpl
veG6tVwT+bsaNscy+HMpIw9FPINjuIB3daaBcxVMXAZlI2kbNhj4YyMMlUU0mTYFOVAjaXxtTX8X
kcXuD4kQT+agHLS6HGBv8KqX+OaOpxUbZ3bA/xj+xSuPd8aa/LPbm09tbO7I0WjGLygG3LcUeBax
JEi6UfQc941N3HJRIOTpOOxuCsOkfqe/I3QQSxdaqs5KCq6lbMveft1bnHC16I1Hu5Q9jQ4TnDRm
h4CzDghE9UMBHDnXnYKdewQZQ+wjeprlTdzpixYLauCpZEE2pBPpG7D3+f7U3bKgH54iqgjw4hWm
ilp2dfbYTc2weHbRzx1YiLht1fd4RDAr58qT/799Ofv3lM+/A0v1goF5j+jbBEvGbpcqFuA/kRx8
OY+Ep00v/SUG0m2+CyOJ/qTrmvFWywv4yWPIMAE5OkxINJN7lpk7zWwpV1kUPK0JWnsMlNetNOwj
Ej9q2rvEy5c1gPYYux0XopDPL9WPM44ysVOEro2/Gk7FFbW0g7xEes38x/pu+cHKgoD8GYret4yk
rWehp+9kco6N0F5QeN9e0tsWtM26/mMuQSmZWDHPMTh0IV51qrs9ZHBDsjSoCaliAsxygRoBY9vz
YYbWr2QaNxDcQ49ZQ6mE+ccmTic4M1XrRbz05eHaQwu4a2NGC8lIqyeSKOdMjXnbA2iLI6EhiEe6
olqGPaaQQFu8hjLAKajOIP0EaHKj8ui6zuv/FVMVpAcp820CCEBeYBzPrARS3P25NcwQ5j0v8tZs
827/Wdhc8f5VmLE7D4jT8zuJ+xGwEYmS6O4U2M+EQ82liiqJq66BH5GDpg9Tq11DpiGG+PIR17wN
mKoYTGj473QHn2OSpU5y4sbKy+rjS4DNH2ue0V4n9Tp41gvICv46XGAVjInoQuvta0CvdkPHT5ET
jTGg/TUiEILoCQbLqb/SomZOpqWiwEdplnz5gcVNv6y0G9/yT3I7/LsGHsNG2c9pVVHWZhmCIPiD
K9q4bEmFo5caw68F9bqByplSe3JOzk7vsHkjjb9ShNGbzuGdaG9cq8MjDFvazPLQo4SoIXUr6Quf
tUnOeWo0VYlCw1jjoK5fO2mzbrCOhGert9NfDTenwTWQZ01hOnZKYiVNFjLoScktYqcWZw0EStf+
gGZoZx6eS69RJpvnLD4JvrrL9JaPJxl+xedCbFeJa2KAWcD48k5q8Wycv59bKpITkob2Qa0JXUn2
DG3rgJf7tfqMuTP6XNH2bemCnMyuDjCchVpGtGZf7x3dJaI+/bv4W2WEkh9MYD2Jl9A9+sNRSfdF
aQJ0cEdAk23b2KaY+K484l37pH3fd+cEui2noJbtx/Pz0T0X6XkFtnPxnTnn2lKtXmkVbUDxYEo3
88RcWVwNTzrIo1WfZga+jad+LCegwnltEaFVh3xf7C7peK5IXmWr4rUunljNTLRJtfimVxZP15nI
p2RkZD+xzzWxJfQRSRYgq9liZN8K8jJYuXkg5bcfknUycRc55PDWDNdXIfoDDLoSXx73lMnLZSbO
aDOyBxcqnvPyO3wX8+IDZMTuE7R747noqSAmZ4dU1rqZDxwiIC7EEodbe/VZx4rVG4vCQN/zw5NW
Tj+GENvbN6Ppt0/G6IWgyR8xrBGrOElRk91LERYPJRlJJbeP5TQ0H1DdVI8PoeO4wO9Z6AzVZGzz
vKMRez9sGEsA7IV4oFu/6SiTbGAtZDAORs8AnUsOK14RmmJsoumdVySbRRtdu8cJ8Q8o0WB8Ks2Z
x/8j8O07k+FoRsrmAaTVXCxR0FWZm5jAiO2n731T+0vmdz48zHtkDiG9Z01ScPsisEMzrbDbJPKC
ole6YdPxmKKJsaDvHr/QhcV9as/7RkL/ScRIZDkS3Sq+wtFVmVcM6azHTxhaRG0eocXbdQBMNqTq
cjxgoqQa8dpRH+hUUWWj+63i2pHEErWrqLsDMlKcqoiczSgEvaFS0ZM3HkKuUyGAzGFYnyjQ0dKG
Lkfe/V9C0/KmSH5YsZ9vLUxU5qmrLoM0ysbIvEA1sxDbK4L6JnNtoWMGYAHVMRjkBLdJ/vBTVpYr
S/IwtJEo1tnzDNhfRHCOWvyCGHgWWb/DrPMfIpP7iNGwV2D9A0PXQQhAXuyA/MROC9DiOkZCVdzL
JyWfojiMGdlk6QgPs81pJEQ2lGP2HakRs1FQKWb4Yc1dSYJfGsr4IUC6M7u1wAe4swCgM6nbNM4Y
Rv8cPGhQFSdVo5jYNNkOdgHEvoUwd1Jq6tGT/SL07c5Jr57j4NE2DvO3nqI2LpQUYbkpwrpDeKil
ZGbKFX3tLb0oqr47GAJjuB9JThPYIbULLGkmwoCJcxOiwywyf2qbhMqlJF4ozZBgwKFuqycCe1Gz
pmAKWraia79AEcHajIrSvAXUKtz+iocIXhOOGleEOvEhJHBwLYCdxP2/J++8cViMSsDADvYrP2+8
QyckWkAx3sGXX+obQyAODMZHHRX/bbkm00BJni5r2feAHbiJ/pc6/HZXjVZeZa+pltOGk+5+G1je
xfoxisT0z1fFHTrkTiKGyG2Ef/3CrMwt0/v4luhb+78qpYsEAkR7KE9IVtDOHsib56Yja+UZwX/o
wHlF4XVxadXJiSbdcit1u4Up+E7TDZpNXyg/WVqj4UtRJpvjGS9v1KU+LlSxJBGWDFmlLsnxgYEh
pCCj5cYkkerLgwxlDTLjHKk1iSHicEJ1zVEVQHQTZ7cIZgX62HWTGGWMgWlF8V0uwu002LC/X8pR
aS0JFBh7cBX6M+KxzZkLRSUq8qF6t80zO+ftFcd0s63n8JI2witEfZCC4i41Eix4JkXQKtlVXm94
9I7kwZrQ9friBnbJP1R06AsOf97o2Aws8At/aJ4sEex3jMTP2nVwOi6Z+Ey/R8ohz4IojV2nYquj
LKw9I7Mr6oPUOjp/d/rBjWyyfb657sYhHnoLwFi5KTbjO+3xlTBPthux92Q0bAtM194wwfvTKwl+
APAEs2YFA+Vgs6rqh2eVX2dHPuEXXezTyXPaDgZoAvcw59M5YwV5Qjarltj1h0EAzKXHrupBQb/H
0dW3S58Qehga04zim1OV31nlnM7HJSLYNnErYAek8WsIN7kPBc2Hs6CC/k1MrwNqhiK5rPCkYTfV
rg9l35qAI3v+brjGia7TItmSkPshcCg3+9S46Gwm+1/rj85xD56sv2QU6tMvsvdPoKPNt6uL8EjW
Gr7i18f0iYe2eotz9ZQX5Z7dwfxfS9ZTdJY5uOTOLqaX7zNotW9P1QhKxMzYO9PvERN/3NdeuGoy
Bq6zT2fdc2dpXmyDGhuPNhh4QBMNhG5xW0XMbSEBH+bkUPlcgM2alb4cZZZ1nmX8i0bJ10M8Qumk
Izx1YgTSLsxrsseJh45PSEgV6y6tvuN5EBh1L2rzWuoWa+T0Oy6oNgcVuCBS7InpA52+Z5rzg2G4
bot29CyGbo6H/eqXswzJmTjBcWKpgXEiTK5eQx2F7MerwZSnBgnE+W7KOHCa3L0wyjG7Tedl2z5p
bbdwo1YYTO+ZMVhH8YTmjrI2iBW6GWmOVxT5Gu1LoY9wQJi3gdVGbHeN5o6SkIYjLbS7ZnQjTrUZ
ePz5f/OcffL0/mBaIBHm+KqqqhGsdV3OW3f6YEsAItdTg/wO5MKCRTapt5OrtlcKCE2/WWVXfFvw
LeRirqM8VZSQ2ZmXJCkuVYdQ7FBrq/BnjJJMl9sSTuhd8OfcUH2TyiZ7OMbobxsuEuOW+/bGihEM
L2Y3qfT261BrwaxJo4pfdOBNQ5aaZINQdSN3bVu4+seEPiNXK6ptwQOPTmgvg+B9kWq0Wd8yrBf+
PiLSRT8EOAXxCiFTT0zgNLUFtf6XH3PjwALPV7NyOHEI9MrffepS1tQSCZmS7/9VUlk5o7icBWVW
Zx96jgKEQEtAyfko725wqzldZ7yXr0yATFguNnzlsixIps54fu59lujSDgzKeJ/IahhJRohQ2r5v
7fMA6DjTeSHa0KSOpOPo1Wwe1x2kYLZQaUCOUvlkU0853OO53YLAl1jKCEnG5DVllkUiuCXoqgoX
gESOuQJ9hDFWKyboAo1+/JNJqwfuLFs+sylNSOWV9mHgH2jHK9ghbkMnamBqrmVnkwZnySE0JvPf
W9vhWTLStRWA2GXvVDlmAUugPOedqYYrfd0flRY/I7IFIlirgP6AonKoXK9PZFKNclNMENgJwv9A
PByzVhrpnd0XCHc7WXnoZSUsVGMH4ncX+7XXpIdN1c9notsHMLCApJYICiQ3Vc1Tb7QeEBn5RhKP
4e61YRMYa67ZJizT8OJy3VBEHgRHiz9v5B6EXokJ0jkDpHJafly5lgdIrgtZvGHdZAl8tVhnlsOV
pU5cHzOP8KqNUvqoIm3DUrJfl4DhEFTrXnxG5vhJZKXKscjrehk3D6g5RpulE9DJ28zBgZ9Xd+px
AQAmwzcrQtdAsOPB2ufAohwXQPbz2MIxl7kDK6cMBDt7guFKkywQkYGjruFSRTk7YCkcqcyv8sPu
/jnHOJFQTD+4gjqCKbo1kBjW04zTcSqOdGKD6fEvycRGLbu9/Vg5WzyOYFsiWyPcZMFFZEvYc/6O
RfxyZh8vRRGlvT+89UNeoV1WUXRof1kUb0PrTCB2nIRiPZosDOyOCQEvLFntNcacOsaQub8iKReu
NynhF2a5RjJCiKDG3FxeyB0h62B50mtILE3kqENat7yEkMeZIkmBlpz8qiYCb9BdywUlhxIutXa7
eWd+l1iNg9X/ikcfH1EhwNREfRnRdEBGKqIu0uxQYzNGcJwpeE5eNgAYTswrKkK1sFfz1J75JWkl
Yb1Pwe6f93J5KnaxHgP5F9hyy0VIv3owDB6yUmjNJw6hQj2WI2Zw7RUX/aykyJas9hc/b/4BiWY0
Ea/VKykrtNopXY5oP2LOntVBeaM+TzYyISf/mrh1M+fFvttMHSVrtNkfWJBagn99nix1SxB+fq91
cXkKLYaiVO4MFRk69os02Rv5ALY3nGzwfzI3NqaptkDu0UdG0LxuW6HyuE7PLHTHO8iX19OKy4D+
rjJ1g7q3ZVSAIsqrZzHGeGR30YFsPHV6iIM0tX00fWac5/WebaKWbdQEhZy7scY/1XlfrsVblUfk
X8zsRHBvu88TkRO/g09VL0XJSk3xs3Y/fSFMJYS8f7DMMIMy+LrSWZHO79jGXedz1FtdSzadREVX
f16GqWCbb5S4sPLSjeIeAltpQJz8M9s4+8dORJL9Y4eCoZHrxpjeP/W5q1Ev7KCA/XmZsiOB7bBd
fYaaSz65ITAmhl93mJUL8ztkfnvGYwc02dYITRigDq2b8EgG1Df7POa5wJGEZOR/QRdqMENoYZip
TgspO7YkQcxahxDEVrhzDacrushBfWEkzwBJBIWGiILA0l9lOu4H2kUSWsAjGkeRdHJJTfEkQYN4
OXelQPAsyEXuTWBYWvdjGwcA4dKafStz5tPnhQHK+BIBsiFw0NpFbZi+iCbMdUMqWLdEEpCY/Y4v
gQYuZRNAsKjDnwJcGlI13TXQWBkiYuB8bCFEC7G/9JYp3wxPTzZYM06VH3P0gVN26+VuoawVR8An
cdo5SD121YmO4xeEwyO5Ega4B204apW3criUL2bo4k2y5W1p2KyqusXDNnnKbV9CgtcL9Pavo08p
OSwkjm3e7lu/DzrC9nGih+K16o9Thc4H7p2z5WE43EbOSB6F1LO3qvkXJvcHX77VQi0V6Lgpw7cu
8uW3AqQgoU/glSNgyewOtuk3v6fo+/c1X9zBIcChsZlA/uBe4Hs3Fuwd1Pk1zDmVbF0X+eSnGmG7
dphBvk1DxQWs2b+DumDq1UhIEXcurGlvitMwYL9hgyiASqwTdy6vhpTI7R8OvdXAZXVewv7AYl4x
P4H44j2yzBSkgjPp0g2Hv+bPJIuTB9pSXoMu8GZifbPh85qZDuCNfvA77wwnQGJgOKlk1/E1rKt9
9aLKYkeQjQAKht0PVFSEipX69Ee01+yyHHK2d++m84J/OdPCwpfT3JomLf/dOpA2iLLAVrb9o5ur
Gm5ZO0QnN6cB37OIXY61EnJ5HaLsYwsMEGIJZ6pZ3w58DsE7o/RAEskXnQCpVW+w0MDnrHdX+5gi
OSUQ63XbhSV64mx6bmLEYO35KpR+q4rzQFKe6N6dH7opXr9EJOUhuLrSGWPvChhnBgglb+THJila
2OcPsldODGHFX3ai+L44MH6BiCWkgxzs5Ef/ILkBjDggf/q5J7nWVrKtxxdFJ7Z6XZQiw7NeFLg7
Un0K9T0Ro9Gmg7dpJ8uI1a2qQWtcMfrtjsPFlkpuMDuTWNHi9xjHFq0XdLiPKu5E+o2ovG8drz5E
oDRCcp8LBzUCe6G/DW25hwIIxXaynryv6ejLLtvvHrJe/0HJsJDzjPV6l/Bz4FOjTL08djux7JpM
WDvHksgEtNac37xt4vyEkhRu3Jhv5ZLus9UVgc9QgMXq6qXCX/YB54tHyfd5WAY5xCufBFIGDvuq
+s+8YfK9P5c10yyFLkKIyrVPMnlR3v88gnarBY767kqyo6baMoGnPyYOWx7I5nNcuU0kTYugZ+IN
i4BHC00tnBGGYNHjdlZSgtBDXe7gEUVnZKM4XNv2+p+P7WZwvQBIwhTsNay0CPuITXmChXbPqJfB
Y87BydeceCuO7Af9KeMhpKtli4tYJp7LS3Dr8S1EuIli8iuN5hyVBgNhsCwQHciETQajYp4qqmjL
viDOXbXGP5tnLxN7gcYkhsfp1zBdfAB71v1I0/x2aEUwJRtRLby5rr+znYvr/BdPuD181mgN4dF5
ta0zxO0Mlwh4f+NiQvU5VHUpxNxnWYbL+5czN+N8rgPD07DXEgDcsVKGqVIOgO99W2/+sX/53iPz
450p3MnKZvUBu69xqsYZAqLXPRHslSqgT45AGIR2jGOmdCI72hXIE1ZppeRhVixBdg62jCqU7gj3
cEGfGTDWQKvdA6sS0Pubab0EBtpw7M6Mt6r6BerwPAf/in5amdllUvY6le71DMDB8CXIzKcgpxvn
PerfbZX1ChTNSzRwUL/nTROadN86URQ7+h/Tj7g19uhUySKwVlpaDgGuxTyDl6RI1K5A4bhRCJAC
IUOhxwhIjZjQCQyouaZPYk7cTS2f40OsYCYkAV8B13zNT6cPF1+Yp4fB+wqWK44U99NiMZmMxwqo
ngARqX6zEYuGUzbrsEhcfPkYdgn33U4SReEnkV1gOf/by1V/WxlkF8yBQQONU04iYbhXZSkRiLDR
aeREG4AbpZKMjmNiYGqimg26RESsRs7tC1ZS0Zy5v6MNllVcyz0czoUmN5jJJtkFtl9LZwhv4B3y
Xtqep4gX6Hukqq/B0paisin/kmM11C0eMKO9V0YAqBfJgzROUrtToRRI7GASg4fJUSnbo9l0ZzlL
ir01mY9G1sXnSvriS3F2lCE4lU2FbZITw+crvYmDrDH4BcRfAkhoDPCxErl9L7d8Ksahl88eSIKb
VbtVm2ogyR0jiPSCez+gZeT+bdNu1FGqtXypwSuadjtiHPsJo3Q1CKMkFvQcOpPphWQmYYGFd197
vIe8Oouihp1zAAn7Dh/Rzz6Dq2ZXxLQBRai68lwFGPd2S/AmRLHKBTSiXh0yo4CVbrO0okcUccFc
hVu/G7oUS/mWW5ZmvrmtFVqNvYasPM8UfeYRMc7w2J2wYS0OWnmvnZOYX1smxZzPMWp0Bx3jTRmY
QoTE3UFdDIp/y0O9+ZVFrZVe+uz4dHOgKR6oeXwiay52ARIBmk0LjOc9QlbHZz7qjr/Pq5jlwMPg
UEWupttvZ0VILDL/DyQYC4mbPUE5DO2rS1na/rPJxBTQlkwGXAF/qeIUqeApMBzo9SkQvHGfM1qx
m8tablqYbo0gPirDPNVZtiQbAAM6FJjR/xBmjuzCOHJ5hjwvZQ9tc3HYtlYcd6g52/SiPJmvpETu
yXqG4DwjUhFFlE1wnu2R7sDaFMsC6MSr6mon/zTzm7Z8khvfm/Or2HFxSweBJt519ps0OGXGid5D
GOrFXBOMQ/j31YXRzDAP0TRlwMTRv2EluP3C+1hKV9AYlgEmqQl3saIdKgGCnO+n/LihRO6izoWO
+DbAM80gSGpj634z6YVHpNVp3opA9q+H01PUdq6Nwd//w3yYb91B4FfGK+FzWRTLDmJCvnZCYDP4
XmtgfX7U9R0mbzOvmUv2nHvcrDgmA/AY2uRRCorreYJ0+69chUY2TxOVBCjgRkhZqQZph9i6bDJa
v5BPv8i1dTmuUpFEEuFNck3hR5FdLw73dBEWkIVm1P2rC+a+s9vsdqaJCXXy0U1+t9lTacmKZReq
Y70qv8SfugpFNQfaDLkYiTTLzsZ008d0FxEkZnI1G9CYCwY7pe6mfIFeIM0jFdL4YUMTLGecf3o4
Gsq5KiXL1dpIiul/oQfpJW7RuMTfRpnBEkwXVLuwKPXzeXyW5QXYJGHPB1XSAxowajqKT0xx2OHj
sI0ofAbzhOZpN7EP7gMVpORgwCGWj50xgcc3EeS55n2K3twSjmwNxNAlix7YWDa2INsdeDS1SR8b
1XOMKLWmk8uJQ65cMHiRgfjJ6VohkVanAhmk8riTGa6j2Bj+A8hQvX4pc0H9odFfEqMsWWuy+xrD
Z7V99dnviSfoExyn32arbiwZj1kWEVFgYsy+4IdgOKu/MH13tSiJm33Yztdz5+mSmA22PudeRs/p
rKsUbLoPDnvz5qoQ6QtLuM0rGp7I4dG0/DuT659b9uJ4sC3u+V620Q+8SusafCirxkaTIi+Qi/xB
dWtIbeOYffzrzl6jnlO3kjcXMWyMVMfMXlUDvJtARe9i4JyUKhxQs6WZphZ4QGXcCcps2GGiJFfs
XriTkV3HlATRLEQt7Nn6yMRXcJapQqHD2Uh2KtS8Sy4MbzyClvqpLaWBi8cSGCRKJfef8d9p9Taf
JrCUTmiwKTMX7QoMBACyzqytQQbGrhn0yLjTns0BRnJIvEhCfP9Bl2wDECxe7TZcLPIqBhaDHh+y
XZ1+/50I+evjJNWmEdla0ob/uMNcCKts/NSGz8z25Qm8rRkoUW70b4gIkIhMaObMmECzRYLq5lPy
KRcZquXD3uUwRI/lLz+P5/UNNqBxdFh6a6TbIytGoITm3o8NrHHk4QKhjy5l/28oOuHEOVHW2JY8
Rb8O7yzdfkTZ+WVmPMkbXf5Mdl2m8ZPMyo+9JIH2Lp8eUkXX59p5NsynnuduNvZEcuUcJp3ZpXo6
sC61UWjPOhAEWFSxXX1ryQk8Qc8BRUodtycSMU3DDc5U8sqlwKW9O5mK/PQB2JptkVWjNRg9eZBm
UiZ/loRjgBsIuzNKw1TkQT82Xl8U2HawUY6eQ0I/qhM6MhLIDtBnh67f8rQwqY1QZwyRRcah+eOK
sbACho8wu7v61gj7yb/XmLBKNBLZx+v5ScFrvMRS44dw3YHaJw72uZKRCTM0MK3ZrzLv+mJY4ezR
J3nyxF5mcPeAyXjMvcYCzH68FJSCaw+Xx7OJAd5FiFaTvHpQYIBI88gPJw3F9b2IVTane2tyZo/G
yQzj5KncR9ZGKhBl/rveySNWSQKp/BEC6DBxGwo55SQipDeCQhYcbXm28vrmqmQR3TFyUjbH+MY8
efLicug9PFVps/HmHetS8RCWPJw+CPSTb/XSkbY5z88cnwM1IbR+gnQ4cxuEfoNFXP4Bf3sTBlQK
LDzy4lVxwsIbHnjWV1rpRW5KOV+32gDpftt9lzIzGj66AkM3fl3iWvtGG+ZqDnD1FooKvtsRniAX
A3VjW3y3qyN49QRSSBrN9XvnaiESciC8AitRskN27SCMTrsQk4UpVeg4zpxWiikOb1RTV7l6igzu
bNWiKnxM9plekpOt66b5CFoDPQmsE0fjWMcuiQhGAmLzzrWsCMGWf1A7vlnJ/N6XtnJtDcH54cZc
uJbhc07MsqRA/Yvah6r+OttCbo4p3ir6F1WT5oCSMpOZ1Vdutc3vbn6yZE6dK1FkiR1gMewn9ORK
xbNGXYGcNMtE+F5agGyw9RuGurefYFXnXPsFwZqrQZO8zxFX/IcoYYEtGgQZZ71ur5+4ATdqZ+vK
3xvqQssjh6tNxj1kzLOpsvh+a/S+H0uerED4esR4VcmFd3x+b2TfwntWPEIF0PJtdk9l0DGiPbID
Td6SMdGK1iTcG3oPQZYpF37fw20+TK/Btef/zBnmDGy8HRnEjqsSj2H5b5oYGW6zEn/WN9nFQrP2
eeE1C0WRCwiQUBjW8WFPNy42YgZ8ZhzLXQSdWpXnRCS6aeB/mDUGNT3oQtDsBtU+SeAZ91dVwsNv
7AA7fyM0Wr++dqT2RK3RWjtr5wfiymPgYSrifV6AVklI9T6Vg55D+roSD4Z9bd56oEuPknFlqEK7
XBsuyqCfqS4ALQCEKR3yUBYD0Ks3sZavoF1yPdh/yKGgSr8cO/4s+TabRxR5PCpZECdc54Ovt0/V
CeIRWmP31Zr6VXu7xGD3bjNZ/hGB0EyAMTmJWsPw2NkXhDvOBTm7V4BxBWV0UC87InmWxYSVQw2L
yG+D0wKXhAfz4T0nrbOuyVuPvpSU26BbYHUsgHCTZgBgQIn01AhV/rExS3zptpkkzHLbYFyQysm3
G+AWVzXMzFD1/sn1qPhp+YgviPHwCYXN0nqYhYHWoSNVSd/TnjnYX+gS7ex380BO+B3Os9kLN/9T
SkSklmvkx59odS5KR/N/7Iu/tpDeMxWpfw5CaAekAkzqZYjQKlnfaOAfTkmNQP8nYsKUBF2IE1+D
/QF0CN7fjJdWE6sgpZDa0TnLn1USqu2LQMTQ8TKt7iLs+1P50fjba9BE4akzTjuuNdXV9W6mvX63
4IXU2Y95Hj82s67Ru8/yKaoJ4W1Ir764emmcrviMScrT7GgcKM18vwJbeJp814FjRiDuGdxZrVJl
C043E2N61s0HQyH6VROI63echzZgEwHl8oVfW/svrilSGtTT+fO8ghKJXRsBnCsfw2hbCJ6YKyKj
LvL/Unog/N69Cg34YZ7UyE/BbV+GtQGW6K2wGRu4t2HMG0XzbPdB9kEMumilSBNEBBZHJIWfR+/S
E8mrziN+L8KNPybqBX6ZK4E9mOo14EhP+qTWzG5YwGtFmhIgFIay0vsH/5H1ifv0KSf5XXlB0R0T
btJ6Z3Bt9syVEkaVQYRvL9cwAb/optUvpOdDdznhLcEYgWwLuVikH5Eo0bNeUmWbRdY4ez0+M7jJ
+DO2gExZKj2mviCiaCmcmEiIxZ4GbBuWstZxCqsF0rlCgOTmmdNIxmO4f1WXrv7kKsNDCjvcwjOT
nw7lkfZBkas0Qmqi9HB5QuUkWTLP9L41HRsEwXs6OQ8Nrp3Si5dTm204
`protect end_protected
