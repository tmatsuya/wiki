`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hksy0AwoxNpXZgHe7l8gadSuz/IC4JAPHSimVYBcXkCK8LEe8iCZWq4LLOrgc79WXipwAYnqj69M
Uf5kLtKmTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g8gasxx4CiwFJicMK6FcOF4v90/vycHQCVuq1gaHhBQ9dqkVU3f05lOsw39GKm8aqw9Xcc96lnPP
qOR2oe4VekCYOLuLS4Mn7CyDtdyESRdt/FeyCKvTL/Glq75Lcn/CkmJu22ffvAmZRSKyyEkh3hEm
+/ZGIX8su0K55k+5fbA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X6ETUAqvIMjJIDWbAmbl1QuSFuOwDyEW8UgSS3T+EnSSfDu+GvhcFVUjQMW5ZY85qoPIkWsdmP5m
COn3eJtJ693ulNg7bqdCLBjyWPTKftqz3tNVIL/PnlHRxd2BlqEUoLKJWnt0NbqM08q0UVQBWLQa
sDPVKOtHW5JL3qzPEd9JBtwU3hilTBZKAw8zjdKLiAjv/rqcKTSXE1Ghw/h4XVO+R+licC/cb8w5
eviacC60HY5lU+CXXyP+R/7yyOxAUGsZA0jdy1N0IBNkdkfOkzNN9Z0bnRZGtLNSvXFZ5+OCrmse
jKouredCITH3nWMI1qoSKUnR6DZo3EE+gkH0ig==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g7onNSps/4WONz9pImy3/1+lstOW//1EGHUnOHWiQJo5yGtWxxf5MzNJCWLcokwcsdM1E8V3EzPX
zf06bbMHxVCw1jQrTw9VJ21e2Rfu3TaYf3LsVheOtY6bWMfqBGcA8egDpvs/krGbLbt+uHy8KsSh
v0yKaNDoOMlDKl8lTrA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QBBOkVVQE6XSganG99o5HX5PTzUuMlGkkAhHUfUk6i0uwWdarazRdietXQjHAkK/iG5cs9R5rOwN
5j6E0kXi3J1OjoyeC61N5KYF07Bu9Xlx45ypTeGMYxMLZCaQK7wHwbCP8jLqw5pZ9JhmQYFXVKwT
nKCWqxIJCCLPlSiYF1BXO3Lc/ztLFl98Bf2mFzhXO2wOzGlmnyMLM0TQpbkhE0NWSWJR+35AJhql
Qov5XHR/6Sn9iDJJwCHWxsPSP3VzT29phgYHhzwI3+lyLFiXq/oXnNZIZoGL3cbIRejpVf23Niuu
JFNhfNDOkYI6BE9r3ku1NsQGPOuKDSwEia9RzQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
vDE86qILrstf0bCEYjiy9yMhvZ60zYHXW7co7MBN6ZpZcGHNdg9Cr+GtR94Ex88b0vlXeTX5EGIh
Tnrt25psRY9fmpg/x1Jafll09TOR4Z07/ySJAugkgvLx4B0Joi9le+4v8qcsjhNTNqppN/0onNcK
cmgcT6zHTabLbIOv5I7KUZFTNtn2Zzi2cGdOP1ceCUHofkXZ9RXajl9ZIYmc2+bfYGnTt1qYNfVC
QkFDTrp7YJof8F2KgrTZws8Jc7K1wibdylFdqlKmhtKida6m5bzeunhuqcrilVZbWpTyWpBz8rRC
zMePWZ4R+46PcKyQoPtwYPVLlcYsBa7zrSAW0WK7Y9ekHHhaV8W71tC2cZT3WS8iKjxhhZRKm/r4
qzUFl6CxyXZ2yZa6cs+wd0+E0Rc+GTF4S5cVmYtbGAu+wKwuCidurN4YO42/xuc++yNTotP3x4jU
FJ90HnokoY6hvOTsDwzlFIHPGMPKpfJRXPeSYLZSNdDih5GOY1vQdlYMQo11ndS5BzCtFoixujMI
WKRn4HEIrnXl3E0oL4txcf6xZkIKslAXI9H2fh+Gw1hHhnTuJ6Q9b6ay3R6/41jusoZuOiR6o5tR
F6GGMKM+O09uF/fqv56LzR+gQoMoH60RU7Jo1wNcCJpsSBqCLoLnumuYOnMkvkIzUElsmkdj5Lmi
BDXMeaOk+ynSVZvScLwene+cfVqUvWl8/nvDtQtvv8PzS8R9VNhlSipKgUQmtJ1H/OuL1m49y5Hc
hy8pFPf6PUzKEgdxFJlXrd/JGEx9zpbrHqOtGnACXWyyS1Sepaea1DP0jbz4X12svIQs4Uco7MiB
mp+/ElfSmeTQiJOQemYn7+hx73BD2BrTcU2ifz3EsyK47AbsbZU3BLSHNt9VsGzsQ003JMqltG/v
Vx+osKu+rwmeOuPgIshg/1a8NmcXip14i1z+LPNimMd0VTySbqvmwOhzyztbHh41hQP9cytu2Irs
ebB4P5NGd0awBoAZpMYtBtamHLWAs+oq/39Qh6piVX5a5YWvdxixnWcUdw2CqdMnwixsV8UjRA4Q
EyAPRZHlp8GuqDwOgy945JDYC5QbX5T9st85iEOh0ZugXlzdy0xIVkJ96qSypSVHa0ixajJiNxB/
a+0kvjduWPFG29OiUTnzYuVaX7MC5ZPJZ9APiI3jRmazI3yJCU3nARQvAUFA9CGJ09l4fCcjlQHh
aTMh1WzzSjYVT9CLZJ8ruunezNaDtX5RHbbq//0F+L2P69YCdQB9u7jhSzLC2yMqsHbKoejqsmiJ
PXbaL0Tz40aAtLly/bT+Rwdcs3UYJBbLHaQMPYHqukNxwMPujkuh0T9Ubs6SdaRIQPuza4PzA+VA
tQJ6c+stosxLtFFHuibCJWJK6qh0G8FDbhnaWDRTMQPVhfvRaWh+5LhFXCLtByFYUegmJQBkG5Fm
KDPkesH2x7+koJSKBZED+kBxJWi5SxCgaDimdDc7tWbJe6knX0o9dnmQ9w0tL+Uj4HNirSUqYyCG
xPbzN+vtTh18sL8erms/pVaCDm2uo7qJHesrUWlbd4Gv7JThMi6XT6lZm3tAk4AEl78xB+nYmp3w
aa5krrnBNmGRlYsLGBdwL2KnGrpBPalmdHQhc7MmQ0l/Poffwy1eIjKWtI9zU2uVVMtw9Z7GCHGX
hUUbwbajUVt0ueu49TflkVxAbwkKgFStla7nNpgfEpZBDjEND8EzPuF3iDePpesJF8LEdnmBmKmy
pVaAhF5KExvKlYLWlg3sq93UH+2XRLSsl/4/EHVaTbdDV7fuocV+gJDW14nS4QizJhXoffiTJl5f
bhuojH/edDJi3MkwWlpNtQugTloYfLmloeZqCzisAHpX6DxO0m83MDc3LjAaMonrnZBWB0s2YavD
JX9uU/4H4h7VnPr6++vV1I0+V6BUlsoBftzhhW1xttWOlG0PXPuHEdexakc0hMzIy73OaoGikhVv
wJnk5U5mPeR+3bTwj+Pzc6u5aJ7OUAxVjai4Bl5EYbk4XqEm3PQ+/IG1lNTjldi9xB1prF60lMdD
0uhnsyUEc7l6oNSIm69JSusQpxHk64ebtDgMatP85Fq+afaKcQa0wqKlIl4etKrbSD5ddQcuWqow
jUFuru6FCaV9veh8CMzQR6s1uOZXBX9We8KIQt+A5xoQrzlTbrL0QwE8t7WqK0WmdkhwI4QVVU75
NLiXwJWHHhNX1bMBCzntlIcT+mDrP2z8taI1s0MOYXXUV+Bu++CtIEAhNys0UbwTZ1Xx87V3+Sqo
G9+O1sKOdEte8lpblekXkPFJdFRrAV7L50fsO6F20pOHERQfTaawEkz5Ox9TljpOiNK3T2Oy3fw8
bhLVYmYqxh5/6rxIWTLgMYMsHQHWLryEfGScDcOwHXVTyYXWKJv8xr+JMPXhhFn1uqdOnX1XuMK1
DJpBxd5oMnsYZejs7ji4kpx/Jwpk25XNi9KGD+S/0cD65jR078Zx33Lyruk2jeouw52ALD7uiGGQ
Dqco9VuSJC0EJSPp8OnNkE2ZUhe+WiRe8+KtfoStdFSDBXVVeDQ9aKMbzcbO14jtH3BA9XHeimnI
aXlW9xEm6llu0PqBQv+81omG9HOYjFsd+tWKhIIh7zXXzY3EqD6tx8VwPUc8SntiR7CT8yrlVuXb
q37Z0I5feKODN9FufrBU0En0SYi2WvK4q7MWRfFVHKJh+dhDjS2CKF7JCiiSsnJASvu5hiEJh/Hv
Qf2XLnytE04+gopF50BAC2GnwIhXMWiSJ1a50lcMCyCscL66QoolNEtbDrQpRQ4torvbKRty4sav
CBDfbMQCWi9lxRFGxP7UHgmK/2F/N2VhkLlV8vNMA+PxPR9QzzeWAKu2WqXjj8bdQSt7/ewF2nHc
KBT2iDX/C2ggBOApgcAhtUuv5UlXRDJN+DMj7e+tAFTh5O/dSp6ErWEOMSWw+dgoBaJBURG7IxKg
vBapiazii27xaIy1RGh5h8Xe6YEzODsIO9dA7VOpet42ni6Tm8m5dh6Top/IjkW8IpKqeBag0O7v
Xn/J/PWktDZiIOqyHqJ16gVxpeXWqOOHQFzM5HQW2ifHuzRAKSWrz+GoWLoINN1nmhNl1MVlQIZN
Z+HIAtZkhqfQOVXXZK6ToKBDLVE5OtJNYvhUvGFnXhf9fR0RKqPnjfRSbbTAqxji+gane9k1aAnp
uHHqG+Ben6v1QW7mEoelG50XQH2Wn+2C3PzV88Kcl4MjHgHisEAoHyWT8t/r0DjNMvZoEQ2mRa50
c6WCXMzfqS2ObzLosrpIxRNe6bx79Xd1z6W23lH8MsWk5opAqs+znBT077IH3a8QccQ2ZiSLvks/
qR6QockN47WgbJFmC/AfoA2Hb3IPimKIxHdg9FsteeFNV/quvf5orAN4C7PLWYOJdd7fLGNPVsjp
BbbocWrtOYDafCOAin67mNu0E1+5e4vcnKiM/OU0SWJhJvlbgK7ahGaUs6xc1olRgpKZrgq4ccp9
JRW9MX5oRV7EhlafvtQxVoXB37cJ9egfq5j03Jl0q5BON2jiuuCCqs3YYVYjIDTtISYiAKVZomFH
U/4LnYw5x+W1r8Os0LqJXObNJJRZzb+wTjNEc0i76bonwM1Q8IoRN3TR5e0K1gVmRLf3v/sz4RB1
oAW/A0QqRKAI/QB1ReiOep8UrcX45wGlDzzS4+owziyhihriCgPL0YJ25gohsHxUANeCR8T0YbVG
USmdi1hEq3PcOd8jZb9AdMf70Y67XQIzsOw7NYw0q7/BWG0f1Tnqf/xyK56MQx7PwcDsNnv7o5mv
F0gkK5XKx2KcGN2bltZxBS1Hup/JFm6E3f1pv4eueto9fiuTMBonIqskSEtWUr3H+8Hd+OYSxd0a
36Ba2kDwkBGgm0XrtIGTmU7i5QX8LxnOFcc/ymrXF+YjXe74aXVQV4t3fK7a81BThzoUT5xDO5fL
CsP55KvGlmxGdvcPOEEIq9kluWIRoS4sOudgd/MmaV+scQmL2uTP+/qWXhAEjto4yiJ5JcdN4SuL
ThAmbY8pSvnImH/Rfulw3fmfvHSgy62wPnauPByUvWxVWrOVSNtQLUWKSc60SJNjlnfbs73c81eQ
a/UHVHKnu518XfmjW4w/5kW5dz/cl+jYLWjU9InlWo/fDY/2xFeP89IQKLjwNhV3qv8/PtAjYvAe
BlTrIXYo2ucgwlTcPp0YIPlK9AELer40Fl5YSeMRDgsxpCrhFTPpoU0n0+otqKAur5PtxhSsIEG2
90qyLNXH3EGnsh1cR52elAKynFlQjOFPopw2p+vQNaZ6QzwjYpKVl40m3bFKjiSxenT1AsfPvvlj
ebTUTGitN6lNoGfsZIv1p0RCRUqxKpldr7phrfvFmuSmCl9XYgtfdf4t28IodzcyuF8n8HBcqvt4
lFd3RxB5MBjIqwYqlOiobAA3luCdAlvlPZIbX5+TRyLkH6OkP5He0VUjGZ1GB4TOGzblbdSIfkWX
pS4W16NeO3Y5Cswp4EMOlphQsi+UtKxOrBwbgJXbwP7SX5Az0akSDfOrps8ZPgM1m0KPPI8JT6WB
mtTm28OiLVbtVtFGernTikVeNCNfRYQSVztZZOsFeM0RomVkwX0CKSPMpTkY589lZW3o5HwmEzng
Sqz+jsvNKtLHFzLXkltDdW/jw2njwiegPvaQMMeMKEtjv4jqgoEi+SXMZHor6vaIpEfIZJWybgiw
iJnHKxknjW2bmMLVMGzk4tSkO6BPa52SN6Y0wg+YxtD061ylEyh2PEYRhGWkjY0ud5YLOI1KwH6A
o4a2p4vVivEr+7aF/nPypwF2KZIXQ5UMTbg+oZT2yWITY8lzbe4xPqrE5nCgR+NYsPj/qIl9sLoO
QPctU5HzTh1RzUG0jbmCjw7XTMGx7/TXnHkqzbUNRFAoE6XRMyIIgnHYQGWpYNPBGzE628eePaG5
y1QuVvhzBhloKgGAoD+4ehc3UotA4JcmnAnVKrKjpb8j5dSmrtqnhsrPaPEimd/AuLJFbSb7+Cjh
pn9CE5VAuyALF8PsMqpROoXzlM89cs+cEZYoTb9V/UHiuwX0kV61b2cjOX3xB0zpdC+XCAP0pC73
EkNisnKUnftf8xXmsyVKdeGzVo/2D17wsb+g6Vf6KI4TXqSDRETBAHfCSe+uCgivXoAQC087P4O5
d371DEqnUeJLAwfSAQPFGIVzWsp9iC/SFn7e8b3J8/zjpX3p3iSXw1LXQYaKaAR/uMbVQjPX0tAq
TE1F9Q9+r87qarecg2m0gBchvrIU3+axgXM1rGRZmluE9+KWsXspGi90F9+cvEITTbUtUiPSELEg
Klq/WFjcbWvYDe2BBiiVLFx4tsYNF5WPf86zWP+osh9OF/R3SFDpaBM6e2P7JgyYrp6IZHIUDpdv
qks3Ua0WceYF7mkF5q0+f2v+xXVvnuUBZ1sPs88iWbfD118ET7w8CgA8lvXTYgPIRfr/nheV5KJF
fHRyP0nr5DDgKhk/ahVVpjGX/8mUUggUtN7jJhSABsPgdMGgf2dg55+QKK4zlNTsVIw2Yh7JUny1
/ryMIo8Kjd11bpvffDVxF4CMDknNYVIJXkuw4saUCTPEJzze9PC46Xo/vV8wKHRMgF70C78370N/
7Sqtlx5/28twseP+rYJ2yJRdWJhO2X4dot+oEiiTkaozgCNCBtP87DVKBdWQ8IA57QluaHc9srvi
+X0SJnXGOlZAmvrIx+twZpTsBdzab8aE2flvorAq8bSljjW4qGqrhRasl3ADR/fcila7wt7P++vW
FrGr4BqjGom9sqo13+OAzAI6SEv/+6COY7a00sOyZTa+RyYZpqIGjTJzrNg4DSoy7Ae1ybA8F1Nt
8PIYjvOkli9go16rmFFtPZ+kZFWbo9iE0rttMI8AuLdRBHQEe5nVaVNiKsBDnTUtflRJv8wba4Xe
1xbLufRn1hJIwRbnG9uvthxY3MpDTddlCNgOB3IQZ24K4dCV7xrO+rX2qEzvRu7dkR31Myf/fLVB
bcLvi7MQEIPRnch/g6X01k3OUo953Y2PpDvCZWhuVdnZGLLcynuOas3hPfhk9Q/A0rbi4YCiLW1X
C4AIP35HivE0YOWfuUpwPcMrB034hG0fPlPzb6bPVzRr9plowvBPiGvn9aanykbbTElxrOmc95UZ
tBOdeZqjBqdaGUt/X8RLeHDQRP1dBB4OMumx6EC4HO25F1OG/IYFdo5lu2lHGaz08phledoYXrUi
wBwKGDCmzko/04m/xjvjhXhT//3sHvvjbibUEoJ8Zyj5H4c/xpQ8zfj03sBVjV4WX2H5YXGJAZ9n
6RD/CQogieybzJpaaUBEGmwQcvcBQae/ROA3K+jt6cirBd65AOVYTKw/E7Ewlbp2cv9UhlJu7cbm
fVSDXwLNWz6HRUXL0oOA3JQyL0HvIJ8uuJZcez5PDw58ZdEDN+voHnWflYC+Y+/4rgwL4kLMuU3m
W87HvdebmmSOY9BMXdxPaoxfM/C3VLq/PFh81CDzY3zXa4P7v/r32gaVQw5yfDSTkJw+HyJ27INJ
xUfZlrhJgEl4VD4EbLAjAmwfrE+dB8Sc32NP+ckcx3yFdFEgW2wGgPx9pJYO2gXc5Hm/iV4lsw1h
X3tv2MTGJ3LWFQNuTN3bDN2VC4v5sPCTQ4kpGhIXpagQrhyJ73Dt0dD5ias6ypoG7/Guhi/mHyVH
6XwU7Ajf1Sxt1jNz75YOWQ6DQCetphVYZcGI5ZAJihBJ3tcaT2HcOSv7ae1IBNDaoR6DR8g4RCUJ
Lc0Uc/+d1O/rmCOZRMDiR6eT56u9ApZw0TRBEy4SSL9KkEr4VGiUHpFXNHxXxlLonNw3QH8TU3Af
ICWBURgc4K67mS5iPhs7yJaRAtIfEEIp0+mmCufAjDwnrUsM+T90NoHPOsdSEqwXXlbpqZAY3Cct
4egX6IiIbBjv23JsB63OePkXOTo5c0DjW76naVN0aJ8QMf7ZeQVTjNgqmXAlobuT8jvAA8gg5IaY
7yHxs2U8rQi1M8rDSEtPmUqhHNBwWm9L49CRH9cLSsnSKYxB1vwt9X5Cnvg46VXVpPkSeuv59KN0
jhF9lP4nsRV6aeNd4LaMJcLGK8pu9EYLG0hgq8UmM4yaRPw0meov1GuF2ABrvMjsgvn/y5fLnzud
IccWZ2sU611qcNEYO5W4AIGf0VLb3Xaj5zKIm2Ng7A7V6UhZENIbfvZ5S+3mKD09XQxFXjTE4FjM
z8x7qi1B5W5+puAsNIHSwBmM+WIjQkS4Q7SES+C2Gnkkl4SgXTZKM9+J9nZoJzMiTXX4LUVd3xJY
/Boi5jkhIqcEq3Sfq7j9BWOCEiqXtSxYwcT2z1TD9oE6Rh2YrkwCFGXn7OtiMC+UWF8356FVDduc
tPtlg7ku8Otku0JuKoVqz3D1SoC0evk+9SpWZobwGm3nGXkAHniuUDSloAkf/shmUWNuOcyiGNZl
7Rs34p+zOdmeS96VkBz9SXdiaHxpRXwVlk/OVBNZ7X7IglL5JxWyfu1qJZYn6MA1QPozmGYNuB0A
DvjwTmov3RsYyvksZKA07CD9eO1G3pBrJ78uCsdFhiAf5WxOiFw2fihzqPPqVMbXVYbPjeLfifWS
S1yjFgNFYwzBGyCUn1WOYqB14UGuY8UTbBLJXeDXtOthRgyUfrg/ISipT5JdM2PapCHJ5yu1me8Y
vOr/ygzQU28F+FC16UM18K/nYEi1sgaYrzEk9ZozKQBvTjDxarDECGY6J4JMmnI6ioPYOTBhcTHz
eybNYLsEs+DauHOclLQPGb8hpqq+BecGQTYvZFkbbIjf/cNkvtVWuhW1qiWWoC++q4/W5ZBqE/65
Jor0Ccgxstbwea/ba1e8kHDkWaCcHN9XqTByd4s2GgLE0Hhbeccc8TLDiycAT13rFJlm0RerINqX
h7R99Wc1+GbAzbbRJQRYhcj5cKrcZK4Btax6VIELKsaPH9/Njyzbk5yCU+ffsBt96wtEM4U80VL+
0vpP0wIuE4FQICtaiXx7HGP9dwFY+iEg0tCoqpMrKgOmhkfMGBt0EoTP0hD1e9IVrXjBMvN3UT/7
3+V+Ejn5eyjXCdyNVEiaEZOEWAqcOPYrxdNUFeqzwHN3jRxwU+ZpwOFYxqVPFXtPcjUrcNGkXW9M
lHGh8+Feq05DdX3ZekMzQUq421SBjqSBn/mx5oDus64NcbSj6xJS8ehkfHQH/zhlwXk17T1LRS9+
USaucJQDEUXcxtirWThwbSiOI5lUnpWJt9r2qXndBEA054ooydzRakzpBhG34E/CtAPRisNGmKzh
44sR9Zki1gIym7yN2l77qz5GT8AOqtibM0ZiJsgCt7VvBf0Cv9xM+CKtu/HZ63VngOyrPP0MPF22
vQkbf5OaegX3Xo4tT+Uy4RA1WxBeDUt5zeuNbjVE5dYMmRM41kVaPwdYB4R1YcpDiwTVzhjb5v0N
3f3AwiHLlB8iaZkHshn7qhqsNS6Q58X6Lly3rW/dImQrwn8qiQ7KgHQyUqKSX9+8UN1kr2bzqBaJ
ltwrLNhmIWBhRQOWepy4DxsKtEJPOt5ujVu+QJi5LTr7QGYEuhQyYhHKCShPAT9v/9GJaBlGTEDi
0/tOnKRGPxkHKTd03vavvJtz0bdHYWOyLMh2Qlm1h58deOHqUmf6tnx1i1YyRh5/lE+Tq+YErLfc
OfWwhfrd9UFLvHq/snfjqdncJKDXFGz2U55OMF4afPEzDjU6vR57qVobgiWq39jq3ch3erTs1DAg
Wat4QEElYCNvsoOLLppM6cOfGdcV44UBCy4kMPqaGLMRE0wWTPrYrhZVloWRERJknOfZ85/DiIPt
65T98Zn7j8abrHnEMPY5wfFguxaU9oyD9D8pz/J7LlPW2X+RJ3i/AJ243W/frww1hx6SZ+3dwekW
UiLjdaKLQ77tFyTAOj2A/DbCq2ln8S4/7HIC8IdnZB2AdGeRgIcK7WxI2zlpjPsVVwwJ0OGoU3Lx
yTLr9Kut3CgwkzmI8BD/h9c8nhDMEvM/JI7n4NqIKpASzkbo5K0Va9cInrJw+gnEx0oC0AisyTzf
IiusQ0ZKfEY3N1IFlmoWAivfe8SOLsVOAdLZ4GwrXlb+d9s8wvZiM8w++1wZkklwshFFWpZuTrri
I6Ukz/rvPjQe5iXlCWUrYunyXbTYW++L8aYYuawvHUZ0nwrfMmbnQ7XBsMIjeawG9yo4JkJSVST6
VHqsT1Ha5t+wA7YJYlyE7Z64+m+A+evj7movbHOeyNiVTxdu1QkNuSi8uw/+LTcSBKoGJvKmQN4l
rBRGxZTK01XLu8VI2Y4N05wNM+XqtBOGIo3CSMCyEd9dfdQ8RRPr1uHnf4/41Az7WXHpf1tGGzh5
s+jp9ECHRPgC3uOW++OlAGUB9ImoK3Ar57R9MhnF/jbP5zHBXT9L3m7ltet6IFiL3kZzODcsSLT8
9fcDnN5NmpP5e/KHa+m/XMGn+V7KyUpLsuRDw9FHsPBnkc2ZZY6OjTScgzjTHZNsSZ9vSfkzubHS
ojyYAaCTyt9SuDNpPuqDTt+Vvqv1AK14HZhUy7j8syUI4UIEfXXHqQ6j4iZI9JWvVc5gsFbaKJke
Yvq6FtNMmw5FtG5PdVi/gEbOjnmP9Bivj8rVxPYp32f4RStbo04z+6kbZm6pOy3ZviIR3CiiG8rL
4hz/u+VA7ZcRIKD9GqL/2Q4pVucabO9RHBIeg55TDDZsaNO3bd6RtqHv/YT78CyiCROrpbaR9ySQ
X3gFRv6fBc18V7ziUOx6qDH12CyaLQ7Tffkzkcyj/9tynBapbSFQy/029hswwDJoZ9IEsdh9wIZH
q426Q6vxqBbhvxDK0kDGatPvonqX3NcXdNkai5AAz+pwk8Jo5wttP+VIw6ZQY/3mSL2qfZBX02Oh
yzmvNKwXLN3r1LI1x+Zc37JwEpj2cThkxc6VV6H6o3o17GDZrkI0aA+72TiX+OqrVq5pBQoeGm6G
upZZI49D7nQDncNFXVclV9ZIsS4RerP0wTTx7z5UMXGfuycs0AS+1z9FIjxQj9FOXDDDdZ8EB7R2
SrwYbWgvGT8RiDXzGR9lQHpaQXfKDWeCOYWL2t+LEnVkzQwOBsFdHb1TtHh5OHC6v+ytNRj/EEuH
sMKdjsecLCkZvAymh6Us3YMI6iB73ees+lyo++S1ip7xlm9ipE0VRM2cBLXhXBz3HkPXEntXzYlg
TNEKE8+rpURv5UKTEZ9bdh3q+gIYq5wwVVbUaEmOIFyb0QTDN/sbPgUm5PwR9Ol/38EvYjHYT4sJ
WiO02wf8QFx2oOYEgMFlWy04H0PnCASpiYbd/ghrCxzOd86PQk906aDwohpPYPP9y6XI7ZzoMP7i
JLEezj2vJDZWHitORgQYXmQCjxDBQvftm3TzffTo+hPZVy2Uh/Dwgh/07OKg+2iKqWJai4eSbvWi
UOqBb0qGP5bkQjKVfrmyuOfPP3DvVBF4ikR6YKzW7O2agENHdHFUPW4ufQrndevlbbH0NRcIrAVr
ZGDx27mO4oKbwz+aOPHgI6+CFZPczm0wbENbegGQ4k40qYS1qRfHZiSWEoQZtLga5E1z5ykw+yD3
/PLoj1qZVrebK2MgJaiYqLbLetYshtP0c44VZbMtqGp2gFgwhxNGvuE04mACCpSjWAyxse3A/RtZ
kXMHr5X1WffHYGcWCf6VbMVmf8Yf35nWf4ZvumS8AkAokY5CXFB1TunZIl2GCSJVWzfjX9gdP/hu
64owuR/lMGGD6OE47cwxUxRyX5VglslngXAw2A8JpVXXNg+m8zTo8rOUL8yb4gxzNP0W0T/cuxHL
0ZFJJkWTbT716C0do2fz3VJQ88B0gBvV0kX9BOrRZORAqq5qanZChjv7bv9db7efCRAG5SsdeMqB
4zjKwsJwjVJKViBB5qcA1q+pKTYSMbNrX6DY0Tx9jeLvyZFEgd8D9Xqxgz501Kb0crvEdWIQXFdF
GVh3iRYm9AqocF01a8RQS8gJ5NVsFRrm0Oh0d3tUut3E9fvd7igdeaIBI2UuNf3MhwNB8yht4t0L
lt5PDVILJo+lNk1d1TOgb8rF08RSBZA1gc9AdGr9ai3si2drj+sCowsEu63KV5BuxpD7zrjSlilW
68u1g6cx2akyNkuW+/2wbNeZ+Da4G281JG6RKnLbPEjsutw3ThNKb07gWI1TsKCuh2aWq+xkzgSh
RBVFhzuKdzJcuJ+Bl2Srmm5rosRZD4XK+5B4+NTDsWycNxkCf69i7gdJ9AJvExHWzCKNSodRNdA2
d//LIBeJql5OWSXAGdvNiDLnJaonOAm24Tx42vq468T0xB1p2PztVtp9nX+kB+ILmW4ZziiDZhJk
k8XzvXYj5+6IhOrB1asukXgL7yO/C19jTPxAkXRL5f6+R7fkXu5y+sCHdaOlpRqzWMX+1jIu61q+
5lYh5RCdkUj0Og+HEUdW5YWJvEOnCVevHPjcZfT36DcWlZAPfhdw4eP5r6Im7mzmdd1RXoRhwiGD
BTW6JFeABSFtB2He3syL/2naXHWCDAFqqvJMtm5B+qJ9WWQlAv0w/oa5KI7Nvd4Izd+gyMKwe2oO
LSgTfmQ6+Zsgd/5JRS28oPIviYgGPvX4kf7QwF8BeoZvY2QDRuKxDsHv9AVohv1hhHnH+qqrKMfA
hVeBGRjszssm0YmvGcpmmiUlZ7/BY9JPxtP1wZmTwleGTS7V2vkT+qxIMyY48e6+x8IUn318+LS6
9ZU8aptawkMUm9T0kmFfndMPleBDG8eGblxanRxBziDR25Y6YP7TBZtfOi5UQTkxx4OAFu/G8ZRH
YZsQ9jljCqZ2pSaV0UQDADAFNpPg6eYy883Kl4Sh6rZ29xGJrSW7MeD0NugLpdO1JnTatDz0dptI
2gs9X1wZZR6tYS+sHqSB1Qm0yGU1OcAQpDhSmOXcYYZC0g0BWuojGlV6WyzOYtv5JBimjEmqHhQi
73+iMXqFigtppIKlBAn2vKKYC3QstEbbaevZLwt/dD0WpPoKsFjosu1RNTqFsR8XEgLlmZngJ/+i
bayvU4X9p5TRSG9mKqocGnOyuLQjv+vxmIjg2taLgd391gUhQ5DXTXBcYYVLgnEdK3a1HtrZAciC
W8p+2joKDP8iaVIriRO7UmuLEQdR0bks4dH+8k1owBD9Lo2/BEj3C64pFCQ92F95s9zA0QBLXyTz
MjT7pFJCG6CiR6Qg3VJlRasSXwkdjJVIiT0KcPYPBelnCHMZPz1Y1NNg9ho+HVbRds1OaAURHT4/
P3H6wbh3pUsXZjtRB6nJulJ8aVwvZMaQ1DV0RPcQzRJtDznkSKg9kHMnX5YAxJrVYLTguzGiAGkV
ezJt67IjBvl+kuStgXatofLfUv57aKdY7D64WCWJizvlGqw30H9dWrox75MgB1BzdhVtkiKTEZ+J
X8AW9HtJWNOBrhCVv9YDfqKDOXMDVt1kBLc7UGL82eJ1Nd4IdkWZmQsLFhm0o7ZVUuqWwZ8GM7Mh
Imlqc2yy7yBmv3vXedBn7QIYIS6Kd98YdyI6Mn9VmUDJpHmgFXg/VDqSknAs57ZKc6yFvSgGyUUc
Fki9pV+3Wi2P7dgQqDI/GAIHCEQfE9jZRDhyl62ywWvW5ZHnA/MqIinCHVu2H/cbiRc0y5ugIU39
t8rpDhGcHKf+lQ0gwjjSO238HIdfbMcuPL4D3yECm4i+OwPcdsQZIwQCVaChb+VyoDeDBw18TqFp
NFssLeHMh+UC0GSL2r7okulKQDH2zm3wDnTWJnAnUfTDajKHdYVnftv1KVObdcbxp/Sagn+MUEYt
RL9GKK5oqxnecT6gRYZY8kmkMrH36F7q9zbHupi1zarQPMAlzrGvGNc4jIlcC2vSOZAi8oT4bH89
NjEDxtHl0950yiA/E5MJsWQk7ne8F30Zjy+SwX8qCMOfnI2MMr8FO3VvqO1ewBkyLVrsrzThrdQX
YaSwRwSAcBjqV7+9kFATdGHm0BX8wpDZTyPwv08+akOEfYlZmHJ0kn+aKQ3MeVobwXYvI8YeBUlG
EjppYHevjMBNXcB5YIW0RfMastNHMg0LBcPIuR7hLPHNgQG27VFJqi4p8KuWNMj9ERuFRG0kblJQ
1udt+UbrHlhkgA6d2ikL2jUGEg3og4Q5FY44JqIsZ9HCyju52/LNV7A67el+czzQD7BQWDcheJr+
P2XZwAwOYFSPQuApeTosCDlhxiCaXjlZ3JjvbdeTsUz4aRMM/COvVDXPIKIzqJDLdNBpGW2EfKHY
Wk2oNsWPlS6LHisC5FmLibjAfB3spKOyUJdGhypz08zg65tkeh7u80XrJsd2P05J4RLOytf0EvNl
luzPJu2MlOh0ChUoZW8MigPJkmp7yrg/2QlN9ns2c8BlLPLc/0LLM5lOx0COZTpXX2y+pqV9p3lV
acoyMDSDQgtTzW03KFe6HuDYOvrG8tX+5y4FCcBhEUHvejs3fSSlu3FSM3ObaifeH3GhwrS2/ZIN
CzG3gwc2TBHT+4sM6VjNpA6hVf8QHdfRV2X+8t3Mu/OGfxlPSMV3A9GYPTm0V/3xOcT7BU8xbT8S
SxUQNHCMDphczAPATiiqccQ1vFGl9GtzlvwlHBNwQLspFhEpj67LhZFQYkQY9zmRMDsZk1gt89Fg
3t+SiOclHtUmruOKBKOXe5lvQwTTpgfIO8VFKFhA0D8AdgAZ4EcYmSzUFSp6avG+YmE6gX8Nn5P4
0kzXOMTyenOQ93nvzmrkR1LVkADHp5kzUkuP2ugJJCktMZYmoeK2WO4Uz5ORBxmFXwOPepm9NZuf
tWQUrEkc653jHv+0daVZLlXLmr4wVuaJUcXl/yAseFeOay6uQdjKpPqS7Rz+HcBStRJHEeSeKJkT
tNtvZC3AReuNNL36MIKPtjEzyBSws/xE3NO8MFwwseIadQq10yDaPDymop7QC18we3zNa3DYAvI7
Hd5IJOmP8fxJpZgjAmjr/6Ej+P60c9mV1xbOgtL30uOM+zqhFuJClwKnV5BqbbVC+OcqCwq4twQA
KEHhjh9b6N0DOCnRnzBR08XS8ciFg5ME4CpkNWJTqgZ1WXUrGmhD17owCi9mjLWIw+1oKnv4ynsi
Wfmrc6/ePMH4EXaeSwYzqrAyMp6bNvHoTEhvKRbhfFbArfgFrNqpT+qifp/jIrVjLe/MLk4hGs0t
MQfurGv7wFdYJIFMdNEy2P/TOJzRcI00xs3m9vmsEHVADM08z2COwovuus0avEZqxdtnJjYxDAFH
6/dB2N8UUfM0Mlz77a6C2Fd6HcPUOa/3NTIMb5MkctzGMhTBRNfc1zOsS91FnJYg6UnD1jpZMQ+T
nQURQ91DoyjHeXpbdVi3FBNpRhf6VHhkG1DcWqdwo3f92lyJ5/PkvD0yA/Uxt3CD1Phi/Xq25ElO
fx25g6ENWFIzrZMzBJTNSoFnN9ah7Fwh7jVNub/rxj0lXuqBSFeqWeXuuY+YoYyUIOaYYXqvHilr
TNtmX67FIXo8XTP5t1KPw4pfCN0CQw9IQW8IZ+5ZGFI+H43jb36j1x12zxnK+iv0XAhDHTxiJLxb
4y9/Co/8gezxJooNnaNpNNocAQhyv6tZj6wdmNorjpjlps2Vcjey92EFdF7cdMlEItqEZVy9DBej
e8aNV8UqDEYodygA7wZERc5djYiwf7Mw7B0/bg9nAqyo7lAN1xt2jjeu3hjNgwDHogGfNJQFBetN
Kcf2XQtL7Q==
`protect end_protected
