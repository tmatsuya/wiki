`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CMnqeZYv+0CptuYfm2JFNTsLOZANWIBjkCPphE0w8DC+J4tf9JEKQRME5gqb6qikKmCeQM7Oh7Jh
16PqsiXOMQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ltiR8ZrKYDBnWuEZKCmjiOcg6wJ6lI/5TAF/9VwF4Q9WVUIK7wAmGhlARiNvQk8cgVef6/rydvh6
CYED+tNk/Wt3kUlwZloUQBVou2+778mVxEhPw80U38ImKbo1EuYqX6koPn9J6W8wYN9dHfAUglt2
7ZB2CbnpTNm496+wBOE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bZ/5epYy7/bc94t2AS4RaBTbp7ND/RRSPj04SPedpGbE/Uo4rPOa6LdL3EijyFPdpgQx8krtERi6
0yHu4qiszTX30Tf9FTYk0HBeDPoRJS81/wmfOhwbe5lYzovgrfFVjhaEpdSnTv5P/nCAXL0CucoE
iG14ylUkOlRV71nQ61YmE4kOYNVC57zxqTIvPautYAaJFqOUGTrCyk+pSSC7RgEPjUYmvYeLtyM8
ZJKD8Qo+Vu11pc6KK7g5a+m/6RYNON9NII3OAvPwKpYffYHHZqJeNKqJli504AfCOg1NnCuRIfbZ
JQty/GygLgQOngznQ5TDwcHfHZA0f9SsRVQMSA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n8g9msMSXZHcqT6wcEvLsP1onUnE5g6Rs+oRelIZzBm29ZGLzAun0xmPRbLnzwnntjWDtTQOf/SL
zWCWtNDuSZfLeM74yvvIXNpnA+z3LQYBDfoP2ABUA8XB4ISy3hUjpWBb/NOvfrrUgjrkspXJQzA9
MbITVr+CjSiJxQ/PnTA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XBNCCqVTQK8eD7Eb5HbrxPqcaLV42qd7O12nbSvVNCmDINRnwsi41RSkPux0hWqmQC2N6TimiAmL
ZM+wk9XX7gbP7uK5/41bfix52HYJkdH/M96l9JvSWRda2uFtEQC0a6S7MJCI8cV2BWIIZdybYEQE
ud3OjqlypR0akZl6GHrJw3GV9DV8/J0e2qvL03DiK55zNlzdn6xyr5x4UYcva8JJQMVTwr2anCGT
eb5VK2bdGou52COHz4XtGWl8DiUr1tbLQMXMf84e1d129IAN+2aeSusmPYxnRKiH4I461TY+e9AB
QSIwL6ZDcktUhksXEytPvQ1ialWOLzjtDbtZgA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15008)
`protect data_block
s2WuA02Y1RBwws6EUqE+HTvfweWK+q0CgA3SZXRG+CptN9BJ3s1RPqVvf2URfU+N3e46KiEjcfDz
vZDel7EFhHKswNrMUOOWfPNrckDnilMcqqnutsoNxy8UqS1lSkxE03MsiApDMnDbJcabS/hb1rEN
CvUlfHbMBQ1UnHQact0gvVogPJCQ19mTOHULC/lN8Nmk+ht1d0b48mKAsFFhfWHobXoru/qNc/Ow
zWRgke5uyjHdWb3n2Z+WYS5Gh2UocU7lVTCNxdxsQfYgLp5LINeszhpWUNNMVRxrm3KJDIK3OoEM
N0G5vxL3ycaaUJH645yX0ALVVzn9wSDfEk//gxHzMDvV3T4vYin/yNPH6exDaQ04tQ+SIX89WC8v
DUemb8U0qXqzfjp9fGM+CNv9yjZi6F6gml0KZI+ZIYgnykR1+kYe3Lszg6RMThs0okt98WHLVNuT
rpo8c2Pk8RH9FkaSg7aJM/i22D7OYCy5xQFXphsvtW/l6jLlKkzRi0xZMuAtFC8OCjHksc+2QXNE
uYPMN2QeWvDF2pTwDgcuT7GpLQ1Iex/Z0Ls77YNlikPJ9mqrMyl5rOORkvLhiVSj/GRfJVXP6wtt
rTrVVl93KDUl+IR4AV2mRjiUSCs6AlQAb5PqE0uEd5krMfkhmwp1I/sIzyM1gps1lfZTaXa3uUb+
1HMHeTb7JVQ+diZOw2LvzEnoO2nBaj4mn7uiudEU5VAJCZAFpUMSG74FatmBmwIhEeHieMpYdH5V
tfxQyN6YtinegRitDCl8/v60OIZHH8GssVWncxpRWBXQ9JjW3ch91oEfyetDSxI1/92Iq+DN4IR6
yP088TwuR6NmFJ1t2aFjKTD2y1rblN+H0MIDslsk1sPX9GPqLwP2zguwxubhUfws9DS/l4GVNcwk
NyuWUBE+o+WFgiDApCJ+qMVXTncdcq0a1NeRmKpeJVOS1hcjxwjMyxFlEhii3SJcBbAd+3D+zZ3o
gIvKICcSOD0mXl8Cb+n0lRmkgNzDE/IosVkg0B3Z5BLCjPvZAcmN5ZEQ9usjJHFz5SRZCK6pPZPG
w3c9rCcPVRDXlPsjT4pugcnGXilxfeUMQy3bE1boGizhvCI14FRVK665I2pTPpTdtLVvfslLmooA
oqFOrF+oaMIHv7piT5ZMYLi6m7WWqmPWJvs9kXWNco6r7v6AYy5BwOt3oCBeCGRdN5KelgZOTEht
MncU5x7WKNYuQASMpmzQxdCRESJUusIRARpWvo0zHIcYFqs9O44F8UDreQOPdyEIvEfzTTWyaeLy
77FYfklRBn/lGvZeCVTHcYnEz9n2HmRu6un0WUcQwsPg68cQaI9fpskxKPho69QGj60oJvpSaIRr
tTPVyKK7nKNoKwLibDufMVhVqVbCWIBkb/X1y30xVgyWqrAxNegMy0yS4teWMOVI/Q6OpdnPTDjH
/RdM9ZDjWUJmmo6YlYqnrtBTfpiNwl1yE9Ws6b9tsCH9HFc/b5EhvBPOPRm3KYdVVrWAOWfHZjeZ
5HbxqzlKwQmmYEYawsmBTns9S8GIuJDmzdpPVym9YzNNcVK9MY1SuMQWZP4GtRlwIEOZT/WoccT6
9hutTooeQBqgjkVJOnDp+BtZl8OJLaZcy2NurgPv14kCpeeqCx2/sP6vKzxpXkKjt386cDxmZzGp
j1moKeicoFokrf9M3mz0JRTZ/G7BnVZ0JYwaSp0kVFQB8EvLPR4kmNNngD3LiMs82dOgNCRwTtQ0
NWUqGX0lEiejmCxW2qrY3N+GCzt/QKmNh5jfAt6rye+5KkZN4iC0vbsdTm886By/W6bfTxH1JC7j
X0rXQTQTrp1TlgfPvBEX4CeycjGLj7YyevJjZmHm1OEaMExzhgl3HQxfHeqhJHqWW34mwvxM1l3p
twxKiLhj4z1J9DYMgrrbxknOZsR7hMr78ywl8e4LMw2givBa9+jH7l9+o4979FbHZvihElorn2zL
qTbfGqFNSC1AZ0r92fgngKB00XK8/sRdOLZQEIWyeQlo+QFmDkGbZG5eNNNGLlBA6QMBEdAuQbDI
Nsu3lv/CsqIedOW866q3zXd0WM/muUs0zAxfX5PqlwLmMK2v9da3M1/u57qiRzSi9TbY2oAvQWQy
YP2RSHEWi6bFV/2lZXiWD1xH3L53QrxCYZ9rrBOMAFPQQb5LCS0eRbz1/PwJNG+YIIU7tUOkbzcI
VdSv2IJQ4Em8Wtq73lfA3HUPyvMXyjMCxG2sNuT9CKENjq3z2vayqsYG8brKLvurvqX8hChQzK2c
nJI7/ftmz0o0O3no4dTkT0tGGCfGoJdcAqy/2NlpG4DIxHroDshy4BeUMR265ccPu9raXKOKjc4L
EgWsLUWRCD72mc/hEh2Qzqowoba6yMYYgZ1XRlFuKqsxJjpU8JX4BuJCNJB3n8aq5sX8MoJlb0JO
VX27R8ojeavokebEb3kTI/4GlwJq6yBxDsOa3awDKoKGyWFqlSsl7QDwhsEIns2yXUQ2q118P6hO
Qqo1Ma9/mc51rRqd3DlhlNRI7mw+7ejcDyYxPgxZpCzMY7Zdx1EAcc5luc501vCYB8izy0w4qpew
msd2Fjjw1AcVljboBA8heyypty3vjvUdEoeUwu1XSycTg7qLmBetTRRUa5lNP7Ng2AX5yxV+jYqh
X7P6bVj8vFNTk9uoPVAIIkSH818bWyym+I0PCcERmp2HC+Bv6dDEk1EAGvMZOgiGgTSgFE/AJDYB
oAWTLKEkp2ZPY6xLc4xaUwFsTtuoIDKkBULpbjJh84BsBgvIoBy11et1YaYIz7detsOwPv/B9oOo
oiTC12nCU7Smp3k3q9vsegxdn1UefM/ENipi8BL+hOwsO/rq0o7ltz3J0uwYnyG1fwC2EayJQiob
0XXqsA8ad0FRVboqFY9FfsLjhJq9eVvJTAQ6oTVXlgOisWA/ohU6ysuDzdzIUOcnPVQeexV2Fddx
BJcAhAIHEn8fvKH0NrK12/4HUWKmzthsmu9kQsFMxcezIxkWn150r+HHC2CyEAj7s+GDXSpOPvLY
3JHamoFjTzlJsCtEFh6G8mSJ6xTstVvl2ydGjeQuD5MifGgcCE7wvJDRk4rcFzLVN6yITi832Ozr
wLzAkX+OmTVr1qh8bsAIWKYWf9jcKrhKFp4zktwwy/mvM8+1HDrCSUkFDpFmbuR61BdGpn4tGeIt
iYWUjKaBiqpiT1I+BBZwtqhRkAh24t+IcMycWrPW3g+49uqgyCNGe50PptOzezU+4XWCu138BKd9
IDogKMiAnVnQygQfONcJf2LwPOIWo4AHgC5xbdYuW8Tq8LST+K5Bty4Ze266Fa1kyFtn0aOyBBOS
m7ZgSaEWZnRz/jDstxJIIuvppPQWgrqveT5Z8qddQ+dk+eTKn2LoNmiKbLU93dGBhwxtllTJSG5i
NVwCaaAsjT7ZCGcQgEsu18vn1e6BSvKVrfJsinbNVUPQ8heWjXUoaocoFYLmDVEeSCrujxSXB5Bz
T5lMNRW+ciwLolYGAXvF1Rd/abBqpOcjdKpG6DvHhRaEZZ0vfph1oBYIb0Uqt/5/7QjWpuMpd7J7
BzIjzwvNN84fiTnRXg8sgXdZP7MnGSs0i90W+FV4scUqvOQFEF0/q1woVViqPml7rywtnl/jiGBG
ca679NAvlFVnkNDc+ggSkzb+0amIdfV81ROEFyZa2vaEQJnUgi8TLC/MZRlqcHQBANLVoP4qjXCE
i+j2YTpPaqi7asfQhpLviSmgV3ZyX208/j/dhOTvrO5nJDXpRqsBrGoJv/+f1mEU2e6vMbX9z/8f
8omjb0vjsdHnWgqBSHWP9vxfwbucqXbD3ujZpy9pbPuBC6vABfwFHnt4FCamciX+3jpOl5yTNIcl
Tw+vIkucaU/MSt78gCY3cKgrxfhRo9ONcyHRnLAmGk3KuKg64FUKZ7n6M4IC56fMjXLePRn5oEFl
e5CxKVTtM5HkHT3eVqBEVyKibqh7klMaSNmMXgdKw4YppT8q/jopeoLcU3Kk1UbZbd4mVAmrD6iW
cC8wOFksj08J5NsYzYfmI07VWKDvaFRUa9hYy3EXdIQQCggbAgrCEQuvCPXVt7xGDKLSoEKNq2tf
F/2vP/vbC7HvmioYErp512v5vh1i0iTRViVQojyxqLY1Uftj9/Ajubhu62EUPV3Wa5cjUvawwBNC
uYBqb9vaPEtn4gTv+jydAUKfLU0mAQLOyhzHpNVtIMIg+MaYjrsdQgwp+AMUh70pulEwNDVna3Wy
IlO1zCo2XSLbdYAp7MdE/ipt3+ddxWXtPf4aWvK12xdLo1Nwy+nwHeEWZ88UoLb7PO5suvdqrlxW
7c6KdF4SnLZ4bHrL2Lq7oRBpXQ9P7cXXZn0kbvrozuoI0K5sV1SRiIFVFEphrNTS+fZsHLfTTyp1
nPPPS84izQOIliEbkUtU8Zq9+NTILs0Z3facy/vRoXu+sysECzi+aqItQ/5hf2DNzmEClX5HjtCV
+1w3Va/4IZ7dvsxkso8H/Y3mqcA2TMRYaRewNnjOjf+G2wpWyJL/bIyreeXdjmZ5BD87vz7HWaAS
0l/vOSlJX/jCMLL5WbIIDuMi3vVIujEqLh2IyGQQrwyIi+KignNVWiTgGspPN9R/2c86yWFrNCNn
DHsb4O1dEXdlbOT/1OFGWbu1mT572tiZwCFSTYOHsBaReWSU+F3nDi/vdhp+Y4032Gs9VcbMwkOK
T4vwdIzUKk22ST8JLOfCuGcquIkzg63leX4W9cJLiGUCMirmyhDgTvgfsUrbIAr5OGWHPHfJSMPX
F83pljXoxF5e9ZSbmKFItjX0jl5hEMQU9U7I1DkVZQkP1roDUPf6K/z8U1Dzi1pDwJmRkAu4zSUf
20p1eiUXV5Jl82VVItQgrZq+8Uy8bsP6qTkcPE9y+mipxiozu9a70USs7clfQq6adA2yIudsUn7l
/493CbdSm+XC7T5M+P0x0d88WBMFOJ6J7QQypQM3E4WGvceRk8v/fdAccIsaVPgmsjPH03EAgWlN
ApeX2mHBPvib06I+ImHYuAOUqNbJ8tgTKVuwK8rNOX6iGEmvTu2uZP8XMy11GrKVbnbQEb5fQHVd
X6gGb2IVlGfXJa22M/TdeLcMLfhTyzjTa9w3eEGCNRVpFDDhBNJpu9yRiFjQPMYxdUiDAuqxsLa5
USJwimgkEWlupVjTBo9+g58Tqivde7ZOmMQ8IPB1xuLtXt8gHIBm5i8Kwyo/SoolyfwugH3aoYhB
C1KfB5DAkkT8xjqPKJhm1uOEniv+bYUXDIKk9PN/Dz+mI14zQoa35KLHRqmVfDxhN10/mKkPDGwz
IBAg0s03rjO8fHe37g8s7qBuuNFmLhFdiwnGL99m75Hr/Oe7UTBxvmslys6eUJKMiWz6FwRS8lbF
eDo132/lyP+S5OuuK7umlMyQOxVKTYYWl8zeBi5RPW9cWEIjyrtYCxnHJW9y15fvHUBskR6c7+CM
d1hIsmIrcy3DnCG6T/TfjQDQM/A3fA/UvzD0bdt1bL+qmgzZ8IltudzApbR+4jY3QRruS2BJ32qP
grLyEYzGQRId7P6XWY3hgbOgE/ph8VBomv5wT8Wtrt1QlCNK45BD1EZ3aKGeGfYMRM9OrGAwET0l
gSDYmXH64BPRQege7N2nJEIdw6V/zOUfWXDBdI67YdVSd6PQyKyRz2Ro78THkn6byfOcyXka2tIu
pPft787H4H9+HKhvb0JInUo3Zq1KvtwhFOrQp3qFnHv+vtFYIVZuUHNa33p6XLoSBxU1zmaXYb63
HsCCCa5tNuYsOA90Ah/lzioMeVyKj4rl2h7nBwrJ62Oo/ymgTqWXKI7jJ/vkBKzugRcCrfaC7SdD
cjzltfMcx5wJPSraXvFWnRId1SRja/SwBFErh5XRhaSkM2er/fKaxS/+fIdZsP0QTVvq+hHpMHrG
CH/FhoT/02NQsALVcWBcbEr97g18NTLC5k0HYjgwxDP/uyt3l6kp5T1+uwS7V3MzyO4X6BowuBID
UcRmDEEdCmyt1eoLJCm/ZJFhko56Z0L9klNySMZjh7ja9IoZOYu2oCIBKMKwJf2ceOWYQ2esYL9O
vo/V1m9nAjXcmbphFrymUPf9LmGsR0Y9ILhCfjHScTh7vS/kl6d7OoE8vTiqmZlIkP+5CAvnchq4
rmevMh4a5bkMGNuAyljDlQCnBLJf7XLmGJSb07XrwvlSsx/MglKbdWcBRCUolF5LIqtJ+tAhC8RF
HiHKeZ3sLtrmmlWxP0979KrIEdCtIttmnUVQS61sKLuqieQu5y1zeGTv/KNHvQh6tHjktzeFGsIf
hWMWZb0FXsPJUsrKRL+ky4lEpbOv2vHdLzq8NPb/umFyNWMrzmRDa5XA+os4VSqkcdLTTEBKQt8v
LK9+xVhVt5KWlRn3jOaxVbfmOaynn9kjNVaOvZHxrartasdf/zvfm2Lru7v8sO90H1f89QJCB2AT
lbpnREV6wQYSpxniqIOWfHQT855iz8UUcnMqUvlyfMUOdJba2krRZb4CJHNYMeYe/3oHTtAPwRPA
u2oUpBGJQhBZAx6lYCPp7KYfl2Ke63h8FgKvPwc9xSLJgcTmqOIVl7dAVXAeBqtf6w005/rvSco1
0HBphXp609oV484+/1ItfK55v/BgdHsEDlbyayPFzbzzDZR4Q3dYFt83TqWGdqfHOHbP9rPUmrQY
2oHnoht1oCLezWFkShE8IRj9zQ7nK4dCYzeefjIIOV+XEdv5Osc/YlQ2nSlJsMS3jmVWgk3jiyyy
4doji5S5UA7jQlFLqqeB9ibdmc8WgU9qzULQlG7J+OKLJQ+AXuvM7TSIXTMrYBK5X+/hsIt5dKUq
Fv56FZAcKcYa9plWpRDe+NfOoc4ZMrRT4EO2LJYwpfkm6RLsQ/kkYi1+c+QuCj01fI/wrhxp1msZ
Ex1fcSH+09eLCw/K4T7wMl+fh3G/gAOdbYuB5Gs4BWislcbMuLc6nP3gTyM0kwbiAeVYeWvPAEuL
+KxA9+/3XGOE8eC2oOs/vML49X9d3P/9CD4uofQ73bBwsUhMMVsR4Pl3YZr9tu8aUNNX2a6+Anrn
iu47gL2uDMi9/5fOSmFEHR5Vhu6ym7wM4cNRnqhSjtL1l7eutqdAKHv+XCv/Y36MXZJwqn6kj0uG
5wDKytPaYezOJZpgtqs56qjE0vIat7BWgPyWkpiHxnTQ1dxDX9XAeP4yqnvoCRPwHNIouJrtj/c+
kRRKOEuhhvg5h8JMigXR1Zvxdqih+dLadni0n1360LIlKihZ6vlZBGDf/KQZStPNAyTs8q1d9vlP
ptWhBXt8NjExf82M5rpaOW5zvx/wgHd925SEiulCtA0JSSTotNm0InfRFFE4YO6v0e0F1PE69M8m
E96JtnkdDQlaKkYaaL9KXDmXLOQFpdBmU/W7x4cLvqd1SWTgiOl/jOOed9ZGXTU8DjxvO06l+kSn
YpLAoYRvfdblBJJmePpNYemz1oiz3B3VUQirtsrfv/SUi2QvHBnMU3Z3Lir3UXPmknpXrqLcXpBh
ehF15pVlH2dplQ1WqvcYXmkp87JEUzIVuAv1uPFAF19rfuSGYX+OM6ruY7IfYJVofDedoeHqY8px
gX+myhU5PvIHCnBP86SuaO2pwMDkgOlGsVdfz54lKI2bmGL+dJ/S4bmqgdZuwsCw16Z24Q91V/a6
i/IVYEDgzzcbPMyHUYfzieNwc6JypAvJTWin1fXm33Gh0y4CzZnYEXKFjDmwfP3nc07USSwZlrjq
ucJTmoMSQthIbPHt+lLvQhWzdkszQGnON+PMACj3IxYJhgGSRC6cw7UwqjCBMYLL8kXsPZpNnnQS
nkeEXoYzqrJHHjyJ86W2TIFeb17RG0amqKmNLyYCxuGixKEn0lEhhvGqhfoJhuSFABkxe3foBn9K
q1TEwCmn1AOb+1RET/oKK6cOljFdHPbH2kQhveQjrBj70fkTEzO5DJUzae0BD7/Iuq7cx7BtAbfo
RSEqpd3SNqagLb8/+k1t4PVZ7BA9UMCviyqEMBVTvTz37PwSFCplZoQK+HwoF596dvsZhuIVwH6A
lLyazzk65UH8orqLVm+Y/11piL8BmYISNIanfVc7y/o7YcX/GBn3/Tsoo+kJwYGSfPELyMMHJRFJ
lMWUsX4PVBASupDW84z2WVlMgzjiY6hayYbc+faSKKCai2/gaZnOYHv2XHtayXdeX+GsH9EOh3B6
q6ln0ya6IE15oA3EILuj9lR0E7ON6AXBNk2LxSYDMi54jucavMcTjiSNxF63UgYxILrNvyvBxOTP
c8v8hNML8GI4yzhJnDJJ9F7bEc9ITdLpPaUOKJsSJzUDQGNd99xMzIzGMJg/fBxSVyaqt1RjYVLo
T5Lh4Z6h/5GbiQK5Cz5JBIBm7mcMoKWHhnOBE2/SlXdFJZo0aozsxcMlU5kJTYm6kryijUqWOxGi
p9B4ICR7nru87FXeptFQzlVPqEzNTATfR/fPrUQmkSA71ST8jfe//dadWxKMahfKnZzcS6E2bn90
bpnN+86/wXRkwODq9KYJFJgQub2Vy+pPoVN/pXJV3oAomjIT8qURFlAtb/s+U6NwI8bqRPd2UTn1
18gtfAD4isBC4QQufW0vPAfq2wCOJbn9NtGwxxLjvoiUp4WvQXE67l2BLGvEw7xRnR+R2nTCbjHD
RHw4SNwR0cSn2ehPsxAhpqiUKEkB+tQ/rLv5p51vdbSgjicFiVSnW8XQDRxxIPzrcdHdS8YJNSDl
cO98cjj3cKMaqK6u5ILCWZx5y78ZLEI0AFrWYq52K3Q00AJl4Ys1Pv74efM43PYqUMr3QJa9UR+C
I0t6pw2uoOiLYEA8mx0/Ogb2rFNMgi3jtaFInYVkS4BNmYmHnfNwDBHLHkcKifwoCumgovP1X3Q0
+0fP1xZK9Q7U0vhFrt9WgnhAiXIe/NIgxVMR5qxonfHq0M3uriUFTLr307ZM/Pc8VCQsvgaQKflq
snqMPTnN4vkKJUpCwzK9nPagdx8+VHRifZseia+V46OiMYt3GDbH2pqaGtji59ltBI1sGzCJDKau
mXUjwB2vNudFPcAIcq99h/ka1mLI6N8Ls5S9Tfz7HY5vdQSlol8y4JfTuk7oiGuQGQCXzkDreHXS
FhWE7sisSRUMtUlwgmEBSFp9vW7dY0epkP9RaW4PlDt6l13Ub4dkQN9bw1XTFkVHH4ilH6GrJ8T1
DGoMgAAL0xfLTU7LuWPrIxS+NlfBynAGAxbKR6KkMqcAqsGZjy8b6cgFiiWcXtENH2FmQMmVP2y8
uYAT5inw6KwhQvzK7gut94/gS83qfMnbYxQ9S8ftyY1CZVgF+JQVoYCN47V2Ril0PZ5HvH3Y66Qv
Dc2ll69HWoRveQObmc0RPMeNyl8yGo1aIlahH6WC42L/ZHEqx89b9es4IIkmWjHj7nVOD60Naw+e
FH1hpYMNkCYhwm6HFaqnW/CzWcswCt8W3Ek5K+XMy9thy0Ko7mbqNCGqY/rZWmwrBkHyg+KVj8wN
NJDOMJs1REITIxWAtqL+l1UWHo8jU+qDSdpWIvqT3iZ6wqvupEDNBjq6PrRtIpmGF2MuaXL7gPdX
yXYQ3LSt6u+uQ6Ohpz/RrqFe/G4TwvIKAVXaZrYqLUR/2t9XBGON2+Qj4/7jjSm8PuNvEcbiEGPr
N0eHuKKbX/WxT+JVAbime+GLqcx3ccl4m2C1Y7yphJanQ1Ttx5BX7zlX9JkcmChX/j/q/JztPf3k
eBZC71CMDrNE+6uE0yZqlyyVrQzgEyjJXtCDNnTqFjFFfIC7UGW4qCKlc3iaGQlMyE9Wg62Xc0Nn
CP31dvtmIKYgeLB85+DzDC8n+S1PvgesktpbmndKWRGyFDHUE4phkOaNC7RIa8C9mghL/dvfZEH5
14w9tB0PNwIM7bGLd7FHuGyE2w1GWxE8llgEfrYA27IvT/jyxzK0xcuKLEM1CLlYxMmtUU5DHFL7
EzAHLjD0zyBj80k1CpTPREGzi7QKhvyEm5XGZu1GXs/czlTrUgK4/T3fh12Rlpz2FUXb2GIahUEN
2RMFSo1A3WFessPs4RBW7DyUghLjoPgJVVxF1NW2hdc4X7XVAlO4K55gpB5Nskl/Av39dM5lOrF4
gMXkhxuo4Ms/K2VbQmJtHGTXzn4ZIcq5yQj8mDfANXcw/4Ud+ATusk5U78kvAKQwqDHdx+6WHA2c
y72V1OTnUoPM6l8EaRKA4nx79TP6sJS/jSdSEtKcwHdwEJi4rV22+mA0DzIo/S8s9aGfETFNZu1f
28E2bpU5aWCL9G8FQJWTr1FDIjikjqv4s3R4iisYLiEYqK/gr2UexBJoPc3I5R97r/RMOWG/l9+5
GlfxWcC4sNljG6zcwoL4DlaUf53IFYZrnwY2g4qF2iWya8vW71GBoj3s8RAcipvWoQkQoL9qSOhL
38w8szdeADBiUny3hBr2TWhzzjG3QjzTgOo8Cztc9JVyyzFCq5Sz9JAGtlad+SqfoRB6Z63FAQrR
VugC/+8AxG6yaZ2V/HYZ458N5uIIceViQIVTMPn2kYeExVHOGmZGZ7Odp/3K0oE5s+WzlDSBGd0w
VPGIgArwdIPcVbzigtn75ftOQOC5y7e4D9snbAYuF7k3SaHxJlTr1j+hJh1Tx6lurfg1UP1Sjyoa
udLb9aCJ1UanH/oyI8rO92w2RLHHnL9JixoGlxJ6gt0excsDkkMTEsRMFeo8RAsaURLG86lOErNM
rl3YqajH/K1PWb1W3Y8quWPHSrKLx6q2KnSAxFTzem3C3YhCtYya8/c+3cQUwTbWP8gcTb+TeJLy
GjlryYweBz+ddCaleSB1pAd1F2/2JOVCdv+EW9YXUBh/h2O186Ikd86Pw9agq+R3Be7NrrG6BBQh
uxTOY31UhOKhofa75HWhSP7DQUa5hdZIpC4793wojX2X8MA/vgPGli5/iJp/F1EB5QJA9Nci8hqg
mDdZbXueXT9F7bPLSb3EjV9FAMICBN1cbiaRG6YhpA8zJcdmi6zpiA4aeorV5sWNRD+W+H/HLBNz
xh4RGR/1xK1tl+4ZORG0Xqine1CWtyNmOOrufESBw+59Mmboqrq1i5GD9IrprehHeqg1J0dw9eZR
RcQQy0DdGbGfH2mGYqiWx6yMa0yCtxovDDxQUyfz196BamFbSgqLAjr4hPjZs45sbns4cwWDw8yC
gW4qlLGQ0J1l54kID9ULTTwBctHXh+bfY1oKU2pY8lBNpXV4mT5SNuiGxXk/aXHoOc6j6iCnwHxT
uByf1ZrleB2QlUkDfftWT7jt5CsJDiQq98Pj+0VLK7z4RQzNOJSkpl/L3gb0TzqrVWQVNfoPaUDq
TyqqTfdrBwT+bnQOYmtubwDZ+ieDuopdqZaOHrkLPDI4UYk1umFOEcT1GpfOM3GJuos98/VhKdfb
TvDz2TgQXJ5I4T1TiJC9JrD/KhV2ace8H5hG7HvoSpWO0kM6ZG/gmDhYwKHl+TmSU9lKaZQtYxxO
0/t506rRcDU5GpsrJ0byCDwwj3xcaClT4VhVIssao2iFhQZuc9nf8rYULMMU+KNfWvn2X1srcN8M
V2u6sSgcC3SBrf3ADzzIbaqOk3kNNSUXL4JhCM4EBNq38KVJVTASBeu3gxB8F/YLDFObNFu0AtAw
TtQb7O+T8cOS6h5hLQSFLQiO4AQkb8hiyWJDEOyFDsSVfhLkpASbuwaLFWvNB7xUKL1A1MdQpHcz
NF8eetT5HGOrL4zlgZ5Q+oNtbwyhSs/ZheUXzwh+8czkfv86epiOIBpX0W/Y6A+/3DkBtKIQu0qE
v0zT4b6JgXWykJ5DrXRDvGEZNuirDdMYUDVamIKlHfPdxSZe+u+C+0mFGPLwhTz11m2eyvt9yDBK
ya1eoWcO3hxyUW+Ytnzm/qUDWWSntX36701SK3d5+96t4tuDo1zo5MCF71mXH5u8w0xbnoyfNt2B
kEoqr0K3nwrfe7grLWXNFaTQneV82j1IjnrI2cqtFOAIyfFEbh/UVgVazzGtKPDuxPWnxw27Lf4R
oySBy4wwkPxdqpvIf5Z01HmnpBQZ+EZFfv7x8JDJhNFv26uqVEuAUVqQBgrtrPwJCASQMiuUUNAx
LzjdTJVnNGCyp+o+FYCj+pT1QqDNj4JaNC8sjlcvzPgFWkA9tJ2hjzii8dTwYfSjyB+/7Dq1ECjF
B3nHM95QQQ7dYVh/wdCiLRrlGnIHckA8bTRIYzW6KTnqXZoBkRGRxcpzJ7s3SglA+Lrc4PM8I+Qb
y6qgpl+bxLyeWNi84vmUzR6kt4wF6vTeSLZpzLSIT3BwQ60UxqobuFN8QYLaUtFASLZgq+2oXWqW
52i4ZvD+oVZ/E7Ooo/g68AHtoRqCFp1HLk4Th45h5cI81EX5w1oVWsPlE+MoLYjJkNMyb77LyUhQ
QxG7GLLqHWwZFc8+p8gkC7E7e3om7LXf8vqyeeFnuDjP9JbR+Sz/HC7p6n3ZjGgz0Hle3E9QEooP
9ZoxsKEsXjAk9heSCarqP9myoBGfdT3HTYUjkU1mMmhJ2sjIuQynuWbs6cSQdoeJf4pKLdj9J9hd
gQ9WfNuP2/+vEyUWuwn2UR9oTfQPW+zBlz7mAjQmzynb5tT4ELTG5NJkPdQZi6w3VdIN4YrwdOnM
V/z4bleer/kB7hKh0ua72TFXO+AwTmYpkBl2lwlhJgrFc+x68Bkj7Z2eVOdDvftnaFEzkTeaJ76a
CHTM7NdIE6hQPBmSMAJBt8klMYoF3h5jY6Ec32uaa+ajDrYHTeTUBNRqPDz79qV5b9i/2rnk6Qek
gPFQhkbrFATAlmTapoDwkYAP362uQU2UuUmi9nQqj3IjHpXY6+BJ7jGV2UiM8K/hDr15Rki7LWy4
49caisSPLg6MgucSW1ClpJxHSdbj+9dbcyIyjwGhCPhPtmubk2hXFvzjrflNjT34wzH+4QnWZ/yL
yicDgOydS9XF7W68oRJyra/0FiMbT2WUEM+LB047zx39/vHyo8WPmdMwJ36bV+sVKk3+PFBTeIYw
ZYqNfV9KNAQI9ctLeOWMD2N0g2WNX50kdusVjwm0a+4cgSFsorFDTie9qitsLl8DGTUdUJpN9ae7
uHpFlzEnJC1N3w0fu+P1OTteCxVj+kyJ35f15ofAdpZVi0TUqv1sBF4GC2gmxWWrVe45XtzwTUoZ
wwhbTG6g3364pln5KVNM2F5vFmDAy9awwnlFWwqvmefFoDz02t3d+QuYQdsxq2sZNvH66AjLaN6j
jdl7EXn7p9U8p5KkVxiiMMbm0IGyDb3rg8CmGj/aiu0jEP9i86mIUoO161gL9yb21msZ5ytnTCtH
qj/9ohmQhko8JrDDJkzMWpupQMSB7myHudXckLqs3DBGnS0Ua0lwsSfM4X0RNzB1TTpQCkDmgK9b
xvSjFNPYNDsfCZH+BObbsL3wC8A7Q4ylMRWOfqilEge4UnmuW3kmVyF4PP4qtimW1VrmBul6sMui
6iV3U2WB7D7pVFkMGSCI6LiJ1qID4UwjyKBU+mLyJxkUo8PZtxtJOchSNPJsJooSFggRWzV6EhZF
1KVXNI+w4yn0RTh165LIOj20i/Wyrv3sCZu+erxJI7PU2RaMKZMq/gEXAc77eJtiMsai3UYmB/JN
sy85gRXaCBuSPLBcarFhhaujJ9txFyZs0uTVhPOX7M4R3RRqS85p/BT1Ab1kQScOxK7F7qbN0T1l
dVJl+dEcCD2LFA6XbDo3MIgzniTIRFZID2/jVWBfH9ZA2T52WGor0Pp1oWyIZOV1HRFpPUgaeZHk
FUeThlXi+9491QllF/0EcIx282hP2MW/gkxJOaJxROpXb7cKdygRvpl4DGkgYHCTrIAW487nBpEE
7E2XkqtQVVEx61WPqFWJbhf8VUs1PAXlo5BFEJfGN5Z0D70YHxS3d5h2OgDHB1q4+lo3N8go48Z8
YiaOw7CVWU9rmGgX+v/b7SR5r0siNjiLSBMcnOzU039j1rMkJ8ILx8s++BEcE+C7+Ch6fmf7Eusu
5ze5l2J9/6SQsEtPgyVWl7sE2xElVQv6vX5LIQvzwEhm+Ptfeebevxdn7hE4c/KnoPuI4QWML+Fb
HsYNrH1TCJXPQgHaSBBFR9jalKsCPqkS27rsgh6DERP0kxQyOKaMbLTbbmzToqJO7NsUeMMDRpWi
MSbK7fPu/dK+ZccuYMbsPbmTAO4DwqYwpyFJHHHvn0U4EAcSeXEJmgApOdjNK9nHQ1AQKd2eZ8mT
CzZUoHkvP0jjm1eQykIY4fxko6RiAGGFNYqC3Pg0Q7dhm1iO/IrwRHnkgIhiqG9mAakASPJv8LQQ
AfFU/8vqrti7UBbPKk2E/HHb5/heBWaEaOaxeW6hcdJJReHFAezErfbLqjemCLn7TGNxsMPLx3xZ
lCtkoMMRZSmL8hhAM19LCR9hRHHhym2SYjWi+2dBmOKBYQlD7688qFBrGqWkv5k+qd9x/a8Trk2e
uGOmJmIKAJpy68Ht8fu08C3mTEYg0Mw3WzmwZ4AyR1/9N+tP4ev5QOa5NCAUeDMLbRZ00iTZC4rK
APE+46rLt16/4bFTl5wlh3uXb4m7k7p9h/Urk6JbJJewNXaqHmLHq7ZJoAMP/MdYC633zs9yAitm
DUMU9nlLtEpfCMIjWJmngNSIoaO9NLOIRbYR6c86wYL8bDGR7eHpw9xqahmUEioEs4Djbx3cpMLd
5/731zXU5u77hFsWDA6nHVKGKzRcsteL89REQVWK2yYHQEOZC9V1XyG5kQYIp17PCUbToY0yvoyS
/WmUKjkoLTOlTvfN9b5rzOhdyQivBUeqYU9fwspaswC+8BacKwObdlSAOSEEzsKQ3J0tfF6Z9Rkf
C+AkTi054Ov2Gj9QxXPovuTiQARs4UYuIXxxd13V0By06n9Fx4wSOaJAplOmgPyP8E1W9oOKT2NL
FEIxbrbAXDeFWBRUf9mvdRyxHXnVerD4yFkGzkBrzsHwUARlNSKyTLVSQo6kyAyTyfMcXz3a7oLM
b3mjM1DWA5ZqAXMZvli0CFmnkO/plxSo9H89lPavjaNSwYmxYBFIIyi1fIWzaltA0srducRDEVrp
XXn99EOD5nsILT8iZpYT5tjxV/oCcjPRjjJ4JfqVAT1zKIEryOmjTtMCFuadyvYCz6Bpev+aNkYH
MW+KuIeiTivkftU9sw3AynFuloeTEOK5hUj/ekiyEsMCapcCCkJq+tJA0vgHsn/mGyjA73OeNf63
f2qC7Vt3aDodV+BI6zk5ccalZbHipOcN3tr2y2i1Tz5BJf5b3nlw8LMfVxVgrLhVW2/hoepfyfys
1VjOuGYtxyA0WnvOGmugcMsRK5bCJH5m0c758mLh2snjcTRnRcX2UCOIQw13K9PBGHi9SIzS5hQ9
r7GHl1rEh0ZpfGt3gRXgXFu6vxaExKjLL9ka1ZwBUOWduMtmLssA/JQMMF/1AIrDTFSWFcsiaVfW
XKRePwjp/89fsjDO+M1vsoRNDn+AOkGzDpd1JIPE+V/ym6i/J8k1e52gbaC9JLiHt9uoli1fvs3R
UOjdzn0qBpMjBylX6QROawx+v4dNQyi5xL4ZNcGNYjhG9f+YVMtlZ7HB04Y7z6ImG+ThOmE0ovIJ
hgX5q6OO3pV7EszZ1BPX/olI5zbb5+ACLPXqEvcPanxXkKJSsMLdLX/UWUt930QAsxnBp3GbgySs
o6nTwAutsWjULs0vE1XTq2uQxaNxfwegz1q1bSqkCU2XVy3rVMGy3YX8w11uOdkz85V69/NdnaTF
Ze2LAG9MaWJJZQF4EqhJcuUNvRe05OKSnO28RZJz5RjFDDCg67zr0a0FzzPKKd2aE14GgYsqk4QZ
6uRtOzvipFiHNcA7adfXvDsr7ySdjIiyPj1GDt8DVMKcQJYQvqmp7xZ3++5wdDXMDT4TTMvu3W2Q
KN8IbXAMHIeoFt/0E6v0kwy23AzxLa/9etCBiZxr0IPfj9WcZhUhS5KcfJUjRTustq3ZOiuhTkJQ
l05EaSqqXoHdWg102cSmVSfEZ/ojoNYhJ2al0KXyv4Vlg4FpNHcgYX3RHSrPyQYJsgXvlJxhpmCB
bYvaN2KJ/hvyVOhPmdG8KPuwoNFAfk091ZCrv9NL/37vNpZKozGU8MYIdhJTTTeHWOi4WMIVkorf
skZyTp7eebaUIoeLbMuyJu3WT6VpTQtGZqwM2F6BgaPlm0LLSP8W7BZhtj55w1ehG62/y6GfP11e
xJKPPf5F08ifBdv4stvIyv3iCAAhZAW4lqVdNi2F5iztwR1n9VpMYx70oXdb1Ftqz/QFNwPm4Xn7
zkJjp7gHUyqYqvu0444lU6shNC+8IC2o6AzPVu0ui91IQkW/6pJuHbST6qK4GatBqz4C+x2i2sDO
kp+M3W7XSJb0j4ur6z4VUMfXISKiaq+hss8fSYUzCd9Ns6wvz+dtNb9SwFFQ9H3qsQrF1tZdg1lm
N7yiFhmj9/2V9G+bTHrUNshDGFGiQlrAuHmzLGaxjgp1eUswZJ7jZMeA95pu5qsRpgIW/GxM3nhN
pBsXM3bMNF0F0sCETVDMl7B98TLC5GwKAUZj76cQRzZvXbwelcRTJFpAoyS0oOZaFKvUdz6X72jx
4lFpbmgSwNQKmbIgB3c+MO3QZMrJEZWUVLkJug9AWoRw/y4JzPzpUzn5uzll2ipSFbolE1u896i2
LgUWnrAAFZB1qaGvEwZ4xsnS6ZO652TCwYFmX872FwwrQYQI+5dVkhEFs4dag0lzP4N/nKIU1Yy1
LPEa0CYr/DXenjvs0vDEcYQbiZX+Yjz489D+GWcJJCKPTgbVEVkm6SnjV9/gQY4JDMOkilzpIuER
+w8TTcKRl0X0WB7/CJySdpJJj74voBo71xHA4VFwdsKt2J09ExymQ4qSuaZpOVIDIweiSucCiaZ3
DHDVuJ1ModHL6/fCSUKDnFKD1jZh1lJMILrmxtJMKAp49s3ExaWdMkwvtx2VCldxteVfoM80DyTP
EzaLcLAzexbgKJcdtGeHSPu//tt1FnGug59sGR8S4iC9+WJ+GGaG0HfyvrugBIlhsAZr5OCVG9Yf
+LQmy7uPPOYHHGKewG/O78zPA5DvWso3CC7sYJxG5qewczR32zl6mkee3kj2+nmsrKPPOpxqBMQF
HSy+3tiXkclZl6acaRyRcXc2YBvXgWJukUjyl1xbvx7uyGHynZ9wZrxF4nHJ83qOoVnjshwAzhXM
yfcyGMv7hAmW3JYFdUQfIkCwYnjH2J+gCTAVW9F3SHGCJBTc4Scemhvo2TL4wiXm0aBSRcjSOqB2
/9ybntVozVOgDpddAm7qR8Y0WSwuHXrk43aBxcKjsZdyXbaXy6RrLoqz53Y1G986Jj2vZ8NfhndS
wEsFeye1YvIrzmM4nYnAsuBg8ioHel10zf/dYmiMtW3gDsKpfektKIL0NyLsd1v4KPXo7IS23l/5
hHk7Bn0SwyPPfqtksM+yp6630gAfgr9M+Djs2FPe23z4QlD1OBLjIC839obi+kLFmbEy5NLUoXIC
VIZmGos0Gaei1AzNs4AIWaP5k9TIfceoF16RQlljpQelzQyR/ja4f/HTmMRsvf2nfJsM3olYbhsS
QZNAJftxLlAwnfPQ6Ofqjyf7IQ9D6ClPieBffdRu3tEsqAs2k5j9dYA7Lup5oyGatAgiLiD08IXl
zNafUPzo/HAphaJrM7oRjErm0r3BgBKbWfRXzSRSg+tUISzft7LP7xT9+BgaSAaKgKaVhxoSEu6w
VzmNTESybpW9NLReLcdjJQHvKS1G+uDgZ2q2mTMmoawGjMHWnzPt8ZkCgmDNuWlyWHUHn9Kha+29
khIyYzQ+55zpCiunlBYKHRELRZXbVCcO07yzkGZWPd9USIIrGXcqd7D09Jk/komv3ZSaSZ9dQ7o+
Yf1jp714fmjB4b0bIz8bFqnlmUHt77F948HMDWL07j7kgluUXjWwrqOAElXE1BglfoRqe0ISvo16
GkJfSl5gpP2u+DMbfbA38JfNti67PO47vI/9WMiAtUkjllkDJi8Ywgb5LDbLVHE/kc8pV5Q5Ns6v
3vH+17lvwbzmZiHGQu517muNQWxoByjDOQTF7mXl8V696pX3Hkyi3Av1jPlVOmdgufaWklH1HTjI
4yAnaVzR0BDY/3txO/4P19eE9BaBX7rHgJ2hZnkoPRBnmZDAIuf5i//BJjgkrdFN217BvpZExOfh
ooRiwIaXLwkY1Ua0GvfCg1elE8x4y7MjJNjiq7sOT1VJU3U8iy2RaX0ko1p6806qDPB7OPmA92sC
RbV1iS9kcg/BOxZ9fv/vrG/HuXj3aoJY8oGcEs5gdxv+eT45nYz6QMjR0yb21alHZTqD4RdUm3Go
gGeGexCyEoZfXh9TYe1HcIi3WdwX/Sr2GdaqHdaZUWgjWsHdlQEtTc0M4OYKUGuvRCyNHql0wPD1
MKpbr9Rz8uy3V608VvoVPWeQWYJ25jGngifqBF6tQnJZHysM0mJYfAFQOffqhHZhgFOjRYQG0vRA
LB0k0TOND3V4N1mrrNuMZIxlRfh1HOsn1KJMZhzds/pmcgYtiJoTPAuySnX/3skwa9jJmeRah9f1
s7weywKrob73QAflabFudHq54Wa7D2cOrJsopFKTh74rpWL4g9A4Mq/VeDA7KbCB5KFIc9uYpQ/2
D9bzQP3Kmq4zBt/W8gdbD1epiAcJ4ZbbXtIWKZ8Cly0vetLPCqaw0YZ6DPZm3jFQEGy1Kmuno7Hc
NbozwXK/xeqtSfpy7hR3OogmajVG8oPH/NGH/ChVQ+IgdbDHiouWBE/MiqjR+7k5Wf1cTH3Db40R
mqeqK+QXHchmlsg6wAEeLxBomt07H0EH3TaGHxgLcQhKy2Jz2/lyYdeEKvew18CFW838iCkv84yV
AhG6PzGuXXEEpU70dX7ctmk+tOmajb9D3D8j092XafwCjaB+p+c+Om8NDQGUUKBs30JTYYoLOgDI
OIZlir4duMMps2VVQ76jM40r1+nV7HbQGaL16GyrjT6rhjlrGcz3dEdjWenWthZehTpO0xGp9vUx
4uOwQIvZskgHsb0UPKeU+hOefTr2gCEhbLbCWAWuQbZlIMJTNPPmnG3NTTsYTPY0pO2boLrvzHXU
6fsOF4U3RUZWOQRMqOsGbOJ1+IEMb/2JTnaH061Kxv5wdV7/8mJTthSwE1GAxJ5AiomavWlV1ql2
AbTamtNHFnzA06trC+Fz6CdqDfyyD4C+jak2ZHm+TBuZq2fHY0DVhOdM8BG0hOYz0WG6XjWXds9g
WGlbnqPcH6rFuXUDZEX1D+pt4YD4uJZItLujN5BrdPdYfqqCR3/wNBV/Kbl+ZxrVvFvZ00IWDwq2
mfTHnLC4p00eCNeXqtfG9BXEJYqN4VUrBAKrNk3lXssHEWcfgr1eGv65Kz2pVZZ5g+HDFSM1Evl7
nO/ZeSJD+KW1woRuO/O4CXeZnPF0P2qPPQIBU5BRZMiNQAx5jM5+puKmLRqV/Y1A7g6xqmX5ZuZC
yhxDc5gjoxu0NzSz1SgIlPmIC+DPnIROhBNsFpxp3lGfPyxdMRjgf5/jUyf4EAy/bvQPQcTi0XH0
WQGwqUKqJdMsjHqX700SFetvwSXHdXZ4MWpZj2ElLAB+sss+lbsem4ncvmRDjP01SxK61ceK4MW2
zrZhg8m635uJkAxwIVmCCcZn1gTIi+Qs9Zj2yXRxTRoU3NfAG9s+2JDK1tXAZN2A4w2S++wkZfPW
hVEbiFZHyZufOrJ2GjTsK9cF5K0OxwajJA+WMWV32kgbKN8U60DHa/ZkoBO7BCf2iO30bkYMLoHf
F3KwZHt3CfE9dfXcnQiUszZoggJ/r4kPi/zF05O/OhkF19HOYMw/guq2JQ1ooi0dQJYwfMvcmlmF
mjoKhkOVWNHEtRLqOd1ZvivdcC9YvM1YqCRGL1vCjOnRK8vqyN5ljvM8mytv7tjGI3fb+tGWZ8PA
A9RYaHbxKcHLPi7NcGC8n/Si/C6Q72WqG0Urb7Ue7itaDzH0oqPqzxcf5eDF6ta9EHt/7r+RfZ6L
AMs07zxmtsjER6hs+GXh+P0=
`protect end_protected
